`timescale 1ns/1ps

module rf ( clk, nrst, rd_addrA, rd_addrB, rd_dataA, rd_dataB, wr_en, wr_addr,
        wr_data );
  input [4:0] rd_addrA;
  input [4:0] rd_addrB;
  output [31:0] rd_dataA;
  output [31:0] rd_dataB;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  input clk, nrst, wr_en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, \r[31][31] ,
         \r[31][30] , \r[31][29] , \r[31][28] , \r[31][27] , \r[31][26] ,
         \r[31][25] , \r[31][24] , \r[31][23] , \r[31][22] , \r[31][21] ,
         \r[31][20] , \r[31][19] , \r[31][18] , \r[31][17] , \r[31][16] ,
         \r[31][15] , \r[31][14] , \r[31][13] , \r[31][12] , \r[31][11] ,
         \r[31][10] , \r[31][9] , \r[31][8] , \r[31][7] , \r[31][6] ,
         \r[31][5] , \r[31][4] , \r[31][3] , \r[31][2] , \r[31][1] ,
         \r[31][0] , \r[30][31] , \r[30][30] , \r[30][29] , \r[30][28] ,
         \r[30][27] , \r[30][26] , \r[30][25] , \r[30][24] , \r[30][23] ,
         \r[30][22] , \r[30][21] , \r[30][20] , \r[30][19] , \r[30][18] ,
         \r[30][17] , \r[30][16] , \r[30][15] , \r[30][14] , \r[30][13] ,
         \r[30][12] , \r[30][11] , \r[30][10] , \r[30][9] , \r[30][8] ,
         \r[30][7] , \r[30][6] , \r[30][5] , \r[30][4] , \r[30][3] ,
         \r[30][2] , \r[30][1] , \r[30][0] , \r[29][31] , \r[29][30] ,
         \r[29][29] , \r[29][28] , \r[29][27] , \r[29][26] , \r[29][25] ,
         \r[29][24] , \r[29][23] , \r[29][22] , \r[29][21] , \r[29][20] ,
         \r[29][19] , \r[29][18] , \r[29][17] , \r[29][16] , \r[29][15] ,
         \r[29][14] , \r[29][13] , \r[29][12] , \r[29][11] , \r[29][10] ,
         \r[29][9] , \r[29][8] , \r[29][7] , \r[29][6] , \r[29][5] ,
         \r[29][4] , \r[29][3] , \r[29][2] , \r[29][1] , \r[29][0] ,
         \r[28][31] , \r[28][30] , \r[28][29] , \r[28][28] , \r[28][27] ,
         \r[28][26] , \r[28][25] , \r[28][24] , \r[28][23] , \r[28][22] ,
         \r[28][21] , \r[28][20] , \r[28][19] , \r[28][18] , \r[28][17] ,
         \r[28][16] , \r[28][15] , \r[28][14] , \r[28][13] , \r[28][12] ,
         \r[28][11] , \r[28][10] , \r[28][9] , \r[28][8] , \r[28][7] ,
         \r[28][6] , \r[28][5] , \r[28][4] , \r[28][3] , \r[28][2] ,
         \r[28][1] , \r[28][0] , \r[27][31] , \r[27][30] , \r[27][29] ,
         \r[27][28] , \r[27][27] , \r[27][26] , \r[27][25] , \r[27][24] ,
         \r[27][23] , \r[27][22] , \r[27][21] , \r[27][20] , \r[27][19] ,
         \r[27][18] , \r[27][17] , \r[27][16] , \r[27][15] , \r[27][14] ,
         \r[27][13] , \r[27][12] , \r[27][11] , \r[27][10] , \r[27][9] ,
         \r[27][8] , \r[27][7] , \r[27][6] , \r[27][5] , \r[27][4] ,
         \r[27][3] , \r[27][2] , \r[27][1] , \r[27][0] , \r[26][31] ,
         \r[26][30] , \r[26][29] , \r[26][28] , \r[26][27] , \r[26][26] ,
         \r[26][25] , \r[26][24] , \r[26][23] , \r[26][22] , \r[26][21] ,
         \r[26][20] , \r[26][19] , \r[26][18] , \r[26][17] , \r[26][16] ,
         \r[26][15] , \r[26][14] , \r[26][13] , \r[26][12] , \r[26][11] ,
         \r[26][10] , \r[26][9] , \r[26][8] , \r[26][7] , \r[26][6] ,
         \r[26][5] , \r[26][4] , \r[26][3] , \r[26][2] , \r[26][1] ,
         \r[26][0] , \r[25][31] , \r[25][30] , \r[25][29] , \r[25][28] ,
         \r[25][27] , \r[25][26] , \r[25][25] , \r[25][24] , \r[25][23] ,
         \r[25][22] , \r[25][21] , \r[25][20] , \r[25][19] , \r[25][18] ,
         \r[25][17] , \r[25][16] , \r[25][15] , \r[25][14] , \r[25][13] ,
         \r[25][12] , \r[25][11] , \r[25][10] , \r[25][9] , \r[25][8] ,
         \r[25][7] , \r[25][6] , \r[25][5] , \r[25][4] , \r[25][3] ,
         \r[25][2] , \r[25][1] , \r[25][0] , \r[24][31] , \r[24][30] ,
         \r[24][29] , \r[24][28] , \r[24][27] , \r[24][26] , \r[24][25] ,
         \r[24][24] , \r[24][23] , \r[24][22] , \r[24][21] , \r[24][20] ,
         \r[24][19] , \r[24][18] , \r[24][17] , \r[24][16] , \r[24][15] ,
         \r[24][14] , \r[24][13] , \r[24][12] , \r[24][11] , \r[24][10] ,
         \r[24][9] , \r[24][8] , \r[24][7] , \r[24][6] , \r[24][5] ,
         \r[24][4] , \r[24][3] , \r[24][2] , \r[24][1] , \r[24][0] ,
         \r[23][31] , \r[23][30] , \r[23][29] , \r[23][28] , \r[23][27] ,
         \r[23][26] , \r[23][25] , \r[23][24] , \r[23][23] , \r[23][22] ,
         \r[23][21] , \r[23][20] , \r[23][19] , \r[23][18] , \r[23][17] ,
         \r[23][16] , \r[23][15] , \r[23][14] , \r[23][13] , \r[23][12] ,
         \r[23][11] , \r[23][10] , \r[23][9] , \r[23][8] , \r[23][7] ,
         \r[23][6] , \r[23][5] , \r[23][4] , \r[23][3] , \r[23][2] ,
         \r[23][1] , \r[23][0] , \r[22][31] , \r[22][30] , \r[22][29] ,
         \r[22][28] , \r[22][27] , \r[22][26] , \r[22][25] , \r[22][24] ,
         \r[22][23] , \r[22][22] , \r[22][21] , \r[22][20] , \r[22][19] ,
         \r[22][18] , \r[22][17] , \r[22][16] , \r[22][15] , \r[22][14] ,
         \r[22][13] , \r[22][12] , \r[22][11] , \r[22][10] , \r[22][9] ,
         \r[22][8] , \r[22][7] , \r[22][6] , \r[22][5] , \r[22][4] ,
         \r[22][3] , \r[22][2] , \r[22][1] , \r[22][0] , \r[21][31] ,
         \r[21][30] , \r[21][29] , \r[21][28] , \r[21][27] , \r[21][26] ,
         \r[21][25] , \r[21][24] , \r[21][23] , \r[21][22] , \r[21][21] ,
         \r[21][20] , \r[21][19] , \r[21][18] , \r[21][17] , \r[21][16] ,
         \r[21][15] , \r[21][14] , \r[21][13] , \r[21][12] , \r[21][11] ,
         \r[21][10] , \r[21][9] , \r[21][8] , \r[21][7] , \r[21][6] ,
         \r[21][5] , \r[21][4] , \r[21][3] , \r[21][2] , \r[21][1] ,
         \r[21][0] , \r[20][31] , \r[20][30] , \r[20][29] , \r[20][28] ,
         \r[20][27] , \r[20][26] , \r[20][25] , \r[20][24] , \r[20][23] ,
         \r[20][22] , \r[20][21] , \r[20][20] , \r[20][19] , \r[20][18] ,
         \r[20][17] , \r[20][16] , \r[20][15] , \r[20][14] , \r[20][13] ,
         \r[20][12] , \r[20][11] , \r[20][10] , \r[20][9] , \r[20][8] ,
         \r[20][7] , \r[20][6] , \r[20][5] , \r[20][4] , \r[20][3] ,
         \r[20][2] , \r[20][1] , \r[20][0] , \r[19][31] , \r[19][30] ,
         \r[19][29] , \r[19][28] , \r[19][27] , \r[19][26] , \r[19][25] ,
         \r[19][24] , \r[19][23] , \r[19][22] , \r[19][21] , \r[19][20] ,
         \r[19][19] , \r[19][18] , \r[19][17] , \r[19][16] , \r[19][15] ,
         \r[19][14] , \r[19][13] , \r[19][12] , \r[19][11] , \r[19][10] ,
         \r[19][9] , \r[19][8] , \r[19][7] , \r[19][6] , \r[19][5] ,
         \r[19][4] , \r[19][3] , \r[19][2] , \r[19][1] , \r[19][0] ,
         \r[18][31] , \r[18][30] , \r[18][29] , \r[18][28] , \r[18][27] ,
         \r[18][26] , \r[18][25] , \r[18][24] , \r[18][23] , \r[18][22] ,
         \r[18][21] , \r[18][20] , \r[18][19] , \r[18][18] , \r[18][17] ,
         \r[18][16] , \r[18][15] , \r[18][14] , \r[18][13] , \r[18][12] ,
         \r[18][11] , \r[18][10] , \r[18][9] , \r[18][8] , \r[18][7] ,
         \r[18][6] , \r[18][5] , \r[18][4] , \r[18][3] , \r[18][2] ,
         \r[18][1] , \r[18][0] , \r[17][31] , \r[17][30] , \r[17][29] ,
         \r[17][28] , \r[17][27] , \r[17][26] , \r[17][25] , \r[17][24] ,
         \r[17][23] , \r[17][22] , \r[17][21] , \r[17][20] , \r[17][19] ,
         \r[17][18] , \r[17][17] , \r[17][16] , \r[17][15] , \r[17][14] ,
         \r[17][13] , \r[17][12] , \r[17][11] , \r[17][10] , \r[17][9] ,
         \r[17][8] , \r[17][7] , \r[17][6] , \r[17][5] , \r[17][4] ,
         \r[17][3] , \r[17][2] , \r[17][1] , \r[17][0] , \r[16][31] ,
         \r[16][30] , \r[16][29] , \r[16][28] , \r[16][27] , \r[16][26] ,
         \r[16][25] , \r[16][24] , \r[16][23] , \r[16][22] , \r[16][21] ,
         \r[16][20] , \r[16][19] , \r[16][18] , \r[16][17] , \r[16][16] ,
         \r[16][15] , \r[16][14] , \r[16][13] , \r[16][12] , \r[16][11] ,
         \r[16][10] , \r[16][9] , \r[16][8] , \r[16][7] , \r[16][6] ,
         \r[16][5] , \r[16][4] , \r[16][3] , \r[16][2] , \r[16][1] ,
         \r[16][0] , \r[15][31] , \r[15][30] , \r[15][29] , \r[15][28] ,
         \r[15][27] , \r[15][26] , \r[15][25] , \r[15][24] , \r[15][23] ,
         \r[15][22] , \r[15][21] , \r[15][20] , \r[15][19] , \r[15][18] ,
         \r[15][17] , \r[15][16] , \r[15][15] , \r[15][14] , \r[15][13] ,
         \r[15][12] , \r[15][11] , \r[15][10] , \r[15][9] , \r[15][8] ,
         \r[15][7] , \r[15][6] , \r[15][5] , \r[15][4] , \r[15][3] ,
         \r[15][2] , \r[15][1] , \r[15][0] , \r[14][31] , \r[14][30] ,
         \r[14][29] , \r[14][28] , \r[14][27] , \r[14][26] , \r[14][25] ,
         \r[14][24] , \r[14][23] , \r[14][22] , \r[14][21] , \r[14][20] ,
         \r[14][19] , \r[14][18] , \r[14][17] , \r[14][16] , \r[14][15] ,
         \r[14][14] , \r[14][13] , \r[14][12] , \r[14][11] , \r[14][10] ,
         \r[14][9] , \r[14][8] , \r[14][7] , \r[14][6] , \r[14][5] ,
         \r[14][4] , \r[14][3] , \r[14][2] , \r[14][1] , \r[14][0] ,
         \r[13][31] , \r[13][30] , \r[13][29] , \r[13][28] , \r[13][27] ,
         \r[13][26] , \r[13][25] , \r[13][24] , \r[13][23] , \r[13][22] ,
         \r[13][21] , \r[13][20] , \r[13][19] , \r[13][18] , \r[13][17] ,
         \r[13][16] , \r[13][15] , \r[13][14] , \r[13][13] , \r[13][12] ,
         \r[13][11] , \r[13][10] , \r[13][9] , \r[13][8] , \r[13][7] ,
         \r[13][6] , \r[13][5] , \r[13][4] , \r[13][3] , \r[13][2] ,
         \r[13][1] , \r[13][0] , \r[12][31] , \r[12][30] , \r[12][29] ,
         \r[12][28] , \r[12][27] , \r[12][26] , \r[12][25] , \r[12][24] ,
         \r[12][23] , \r[12][22] , \r[12][21] , \r[12][20] , \r[12][19] ,
         \r[12][18] , \r[12][17] , \r[12][16] , \r[12][15] , \r[12][14] ,
         \r[12][13] , \r[12][12] , \r[12][11] , \r[12][10] , \r[12][9] ,
         \r[12][8] , \r[12][7] , \r[12][6] , \r[12][5] , \r[12][4] ,
         \r[12][3] , \r[12][2] , \r[12][1] , \r[12][0] , \r[11][31] ,
         \r[11][30] , \r[11][29] , \r[11][28] , \r[11][27] , \r[11][26] ,
         \r[11][25] , \r[11][24] , \r[11][23] , \r[11][22] , \r[11][21] ,
         \r[11][20] , \r[11][19] , \r[11][18] , \r[11][17] , \r[11][16] ,
         \r[11][15] , \r[11][14] , \r[11][13] , \r[11][12] , \r[11][11] ,
         \r[11][10] , \r[11][9] , \r[11][8] , \r[11][7] , \r[11][6] ,
         \r[11][5] , \r[11][4] , \r[11][3] , \r[11][2] , \r[11][1] ,
         \r[11][0] , \r[10][31] , \r[10][30] , \r[10][29] , \r[10][28] ,
         \r[10][27] , \r[10][26] , \r[10][25] , \r[10][24] , \r[10][23] ,
         \r[10][22] , \r[10][21] , \r[10][20] , \r[10][19] , \r[10][18] ,
         \r[10][17] , \r[10][16] , \r[10][15] , \r[10][14] , \r[10][13] ,
         \r[10][12] , \r[10][11] , \r[10][10] , \r[10][9] , \r[10][8] ,
         \r[10][7] , \r[10][6] , \r[10][5] , \r[10][4] , \r[10][3] ,
         \r[10][2] , \r[10][1] , \r[10][0] , \r[9][31] , \r[9][30] ,
         \r[9][29] , \r[9][28] , \r[9][27] , \r[9][26] , \r[9][25] ,
         \r[9][24] , \r[9][23] , \r[9][22] , \r[9][21] , \r[9][20] ,
         \r[9][19] , \r[9][18] , \r[9][17] , \r[9][16] , \r[9][15] ,
         \r[9][14] , \r[9][13] , \r[9][12] , \r[9][11] , \r[9][10] , \r[9][9] ,
         \r[9][8] , \r[9][7] , \r[9][6] , \r[9][5] , \r[9][4] , \r[9][3] ,
         \r[9][2] , \r[9][1] , \r[9][0] , \r[8][31] , \r[8][30] , \r[8][29] ,
         \r[8][28] , \r[8][27] , \r[8][26] , \r[8][25] , \r[8][24] ,
         \r[8][23] , \r[8][22] , \r[8][21] , \r[8][20] , \r[8][19] ,
         \r[8][18] , \r[8][17] , \r[8][16] , \r[8][15] , \r[8][14] ,
         \r[8][13] , \r[8][12] , \r[8][11] , \r[8][10] , \r[8][9] , \r[8][8] ,
         \r[8][7] , \r[8][6] , \r[8][5] , \r[8][4] , \r[8][3] , \r[8][2] ,
         \r[8][1] , \r[8][0] , \r[7][31] , \r[7][30] , \r[7][29] , \r[7][28] ,
         \r[7][27] , \r[7][26] , \r[7][25] , \r[7][24] , \r[7][23] ,
         \r[7][22] , \r[7][21] , \r[7][20] , \r[7][19] , \r[7][18] ,
         \r[7][17] , \r[7][16] , \r[7][15] , \r[7][14] , \r[7][13] ,
         \r[7][12] , \r[7][11] , \r[7][10] , \r[7][9] , \r[7][8] , \r[7][7] ,
         \r[7][6] , \r[7][5] , \r[7][4] , \r[7][3] , \r[7][2] , \r[7][1] ,
         \r[7][0] , \r[6][31] , \r[6][30] , \r[6][29] , \r[6][28] , \r[6][27] ,
         \r[6][26] , \r[6][25] , \r[6][24] , \r[6][23] , \r[6][22] ,
         \r[6][21] , \r[6][20] , \r[6][19] , \r[6][18] , \r[6][17] ,
         \r[6][16] , \r[6][15] , \r[6][14] , \r[6][13] , \r[6][12] ,
         \r[6][11] , \r[6][10] , \r[6][9] , \r[6][8] , \r[6][7] , \r[6][6] ,
         \r[6][5] , \r[6][4] , \r[6][3] , \r[6][2] , \r[6][1] , \r[6][0] ,
         \r[5][31] , \r[5][30] , \r[5][29] , \r[5][28] , \r[5][27] ,
         \r[5][26] , \r[5][25] , \r[5][24] , \r[5][23] , \r[5][22] ,
         \r[5][21] , \r[5][20] , \r[5][19] , \r[5][18] , \r[5][17] ,
         \r[5][16] , \r[5][15] , \r[5][14] , \r[5][13] , \r[5][12] ,
         \r[5][11] , \r[5][10] , \r[5][9] , \r[5][8] , \r[5][7] , \r[5][6] ,
         \r[5][5] , \r[5][4] , \r[5][3] , \r[5][2] , \r[5][1] , \r[5][0] ,
         \r[4][31] , \r[4][30] , \r[4][29] , \r[4][28] , \r[4][27] ,
         \r[4][26] , \r[4][25] , \r[4][24] , \r[4][23] , \r[4][22] ,
         \r[4][21] , \r[4][20] , \r[4][19] , \r[4][18] , \r[4][17] ,
         \r[4][16] , \r[4][15] , \r[4][14] , \r[4][13] , \r[4][12] ,
         \r[4][11] , \r[4][10] , \r[4][9] , \r[4][8] , \r[4][7] , \r[4][6] ,
         \r[4][5] , \r[4][4] , \r[4][3] , \r[4][2] , \r[4][1] , \r[4][0] ,
         \r[3][31] , \r[3][30] , \r[3][29] , \r[3][28] , \r[3][27] ,
         \r[3][26] , \r[3][25] , \r[3][24] , \r[3][23] , \r[3][22] ,
         \r[3][21] , \r[3][20] , \r[3][19] , \r[3][18] , \r[3][17] ,
         \r[3][16] , \r[3][15] , \r[3][14] , \r[3][13] , \r[3][12] ,
         \r[3][11] , \r[3][10] , \r[3][9] , \r[3][8] , \r[3][7] , \r[3][6] ,
         \r[3][5] , \r[3][4] , \r[3][3] , \r[3][2] , \r[3][1] , \r[3][0] ,
         \r[2][31] , \r[2][30] , \r[2][29] , \r[2][28] , \r[2][27] ,
         \r[2][26] , \r[2][25] , \r[2][24] , \r[2][23] , \r[2][22] ,
         \r[2][21] , \r[2][20] , \r[2][19] , \r[2][18] , \r[2][17] ,
         \r[2][16] , \r[2][15] , \r[2][14] , \r[2][13] , \r[2][12] ,
         \r[2][11] , \r[2][10] , \r[2][9] , \r[2][8] , \r[2][7] , \r[2][6] ,
         \r[2][5] , \r[2][4] , \r[2][3] , \r[2][2] , \r[2][1] , \r[2][0] ,
         \r[1][31] , \r[1][30] , \r[1][29] , \r[1][28] , \r[1][27] ,
         \r[1][26] , \r[1][25] , \r[1][24] , \r[1][23] , \r[1][22] ,
         \r[1][21] , \r[1][20] , \r[1][19] , \r[1][18] , \r[1][17] ,
         \r[1][16] , \r[1][15] , \r[1][14] , \r[1][13] , \r[1][12] ,
         \r[1][11] , \r[1][10] , \r[1][9] , \r[1][8] , \r[1][7] , \r[1][6] ,
         \r[1][5] , \r[1][4] , \r[1][3] , \r[1][2] , \r[1][1] , \r[1][0] , n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303;
  assign N11 = rd_addrA[0];
  assign N12 = rd_addrA[1];
  assign N13 = rd_addrA[2];
  assign N14 = rd_addrA[3];
  assign N15 = rd_addrA[4];
  assign N16 = rd_addrB[0];
  assign N17 = rd_addrB[1];
  assign N18 = rd_addrB[2];
  assign N19 = rd_addrB[3];
  assign N20 = rd_addrB[4];

  DFFARX1 \r_reg[31][31]  ( .D(n1071), .CLK(clk), .RSTB(n2211), .Q(\r[31][31] ) );
  DFFARX1 \r_reg[31][30]  ( .D(n1070), .CLK(clk), .RSTB(n2211), .Q(\r[31][30] ) );
  DFFARX1 \r_reg[31][29]  ( .D(n1069), .CLK(clk), .RSTB(n2211), .Q(\r[31][29] ) );
  DFFARX1 \r_reg[31][28]  ( .D(n1068), .CLK(clk), .RSTB(n2211), .Q(\r[31][28] ) );
  DFFARX1 \r_reg[31][27]  ( .D(n1067), .CLK(clk), .RSTB(n2211), .Q(\r[31][27] ) );
  DFFARX1 \r_reg[31][26]  ( .D(n1066), .CLK(clk), .RSTB(n2211), .Q(\r[31][26] ) );
  DFFARX1 \r_reg[31][25]  ( .D(n1065), .CLK(clk), .RSTB(n2211), .Q(\r[31][25] ) );
  DFFARX1 \r_reg[31][24]  ( .D(n1064), .CLK(clk), .RSTB(n2211), .Q(\r[31][24] ) );
  DFFARX1 \r_reg[31][23]  ( .D(n1063), .CLK(clk), .RSTB(n2211), .Q(\r[31][23] ) );
  DFFARX1 \r_reg[31][22]  ( .D(n1062), .CLK(clk), .RSTB(n2211), .Q(\r[31][22] ) );
  DFFARX1 \r_reg[31][21]  ( .D(n1061), .CLK(clk), .RSTB(n2211), .Q(\r[31][21] ) );
  DFFARX1 \r_reg[31][20]  ( .D(n1060), .CLK(clk), .RSTB(n2211), .Q(\r[31][20] ) );
  DFFARX1 \r_reg[31][19]  ( .D(n1059), .CLK(clk), .RSTB(n2212), .Q(\r[31][19] ) );
  DFFARX1 \r_reg[31][18]  ( .D(n1058), .CLK(clk), .RSTB(n2212), .Q(\r[31][18] ) );
  DFFARX1 \r_reg[31][17]  ( .D(n1057), .CLK(clk), .RSTB(n2212), .Q(\r[31][17] ) );
  DFFARX1 \r_reg[31][16]  ( .D(n1056), .CLK(clk), .RSTB(n2212), .Q(\r[31][16] ) );
  DFFARX1 \r_reg[31][15]  ( .D(n1055), .CLK(clk), .RSTB(n2212), .Q(\r[31][15] ) );
  DFFARX1 \r_reg[31][14]  ( .D(n1054), .CLK(clk), .RSTB(n2212), .Q(\r[31][14] ) );
  DFFARX1 \r_reg[31][13]  ( .D(n1053), .CLK(clk), .RSTB(n2212), .Q(\r[31][13] ) );
  DFFARX1 \r_reg[31][12]  ( .D(n1052), .CLK(clk), .RSTB(n2212), .Q(\r[31][12] ) );
  DFFARX1 \r_reg[31][11]  ( .D(n1051), .CLK(clk), .RSTB(n2212), .Q(\r[31][11] ) );
  DFFARX1 \r_reg[31][10]  ( .D(n1050), .CLK(clk), .RSTB(n2212), .Q(\r[31][10] ) );
  DFFARX1 \r_reg[31][9]  ( .D(n1049), .CLK(clk), .RSTB(n2212), .Q(\r[31][9] )
         );
  DFFARX1 \r_reg[31][8]  ( .D(n1048), .CLK(clk), .RSTB(n2212), .Q(\r[31][8] )
         );
  DFFARX1 \r_reg[31][7]  ( .D(n1047), .CLK(clk), .RSTB(n2213), .Q(\r[31][7] )
         );
  DFFARX1 \r_reg[31][6]  ( .D(n1046), .CLK(clk), .RSTB(n2213), .Q(\r[31][6] )
         );
  DFFARX1 \r_reg[31][5]  ( .D(n1045), .CLK(clk), .RSTB(n2213), .Q(\r[31][5] )
         );
  DFFARX1 \r_reg[31][4]  ( .D(n1044), .CLK(clk), .RSTB(n2213), .Q(\r[31][4] )
         );
  DFFARX1 \r_reg[31][3]  ( .D(n1043), .CLK(clk), .RSTB(n2213), .Q(\r[31][3] )
         );
  DFFARX1 \r_reg[31][2]  ( .D(n1042), .CLK(clk), .RSTB(n2213), .Q(\r[31][2] )
         );
  DFFARX1 \r_reg[31][1]  ( .D(n1041), .CLK(clk), .RSTB(n2213), .Q(\r[31][1] )
         );
  DFFARX1 \r_reg[31][0]  ( .D(n1040), .CLK(clk), .RSTB(n2213), .Q(\r[31][0] )
         );
  DFFARX1 \r_reg[30][31]  ( .D(n1039), .CLK(clk), .RSTB(n2213), .Q(\r[30][31] ) );
  DFFARX1 \r_reg[30][30]  ( .D(n1038), .CLK(clk), .RSTB(n2213), .Q(\r[30][30] ) );
  DFFARX1 \r_reg[30][29]  ( .D(n1037), .CLK(clk), .RSTB(n2213), .Q(\r[30][29] ) );
  DFFARX1 \r_reg[30][28]  ( .D(n1036), .CLK(clk), .RSTB(n2213), .Q(\r[30][28] ) );
  DFFARX1 \r_reg[30][27]  ( .D(n1035), .CLK(clk), .RSTB(n2214), .Q(\r[30][27] ) );
  DFFARX1 \r_reg[30][26]  ( .D(n1034), .CLK(clk), .RSTB(n2214), .Q(\r[30][26] ) );
  DFFARX1 \r_reg[30][25]  ( .D(n1033), .CLK(clk), .RSTB(n2214), .Q(\r[30][25] ) );
  DFFARX1 \r_reg[30][24]  ( .D(n1032), .CLK(clk), .RSTB(n2214), .Q(\r[30][24] ) );
  DFFARX1 \r_reg[30][23]  ( .D(n1031), .CLK(clk), .RSTB(n2214), .Q(\r[30][23] ) );
  DFFARX1 \r_reg[30][22]  ( .D(n1030), .CLK(clk), .RSTB(n2214), .Q(\r[30][22] ) );
  DFFARX1 \r_reg[30][21]  ( .D(n1029), .CLK(clk), .RSTB(n2214), .Q(\r[30][21] ) );
  DFFARX1 \r_reg[30][20]  ( .D(n1028), .CLK(clk), .RSTB(n2214), .Q(\r[30][20] ) );
  DFFARX1 \r_reg[30][19]  ( .D(n1027), .CLK(clk), .RSTB(n2214), .Q(\r[30][19] ) );
  DFFARX1 \r_reg[30][18]  ( .D(n1026), .CLK(clk), .RSTB(n2214), .Q(\r[30][18] ) );
  DFFARX1 \r_reg[30][17]  ( .D(n1025), .CLK(clk), .RSTB(n2214), .Q(\r[30][17] ) );
  DFFARX1 \r_reg[30][16]  ( .D(n1024), .CLK(clk), .RSTB(n2214), .Q(\r[30][16] ) );
  DFFARX1 \r_reg[30][15]  ( .D(n1023), .CLK(clk), .RSTB(n2215), .Q(\r[30][15] ) );
  DFFARX1 \r_reg[30][14]  ( .D(n1022), .CLK(clk), .RSTB(n2215), .Q(\r[30][14] ) );
  DFFARX1 \r_reg[30][13]  ( .D(n1021), .CLK(clk), .RSTB(n2215), .Q(\r[30][13] ) );
  DFFARX1 \r_reg[30][12]  ( .D(n1020), .CLK(clk), .RSTB(n2215), .Q(\r[30][12] ) );
  DFFARX1 \r_reg[30][11]  ( .D(n1019), .CLK(clk), .RSTB(n2215), .Q(\r[30][11] ) );
  DFFARX1 \r_reg[30][10]  ( .D(n1018), .CLK(clk), .RSTB(n2215), .Q(\r[30][10] ) );
  DFFARX1 \r_reg[30][9]  ( .D(n1017), .CLK(clk), .RSTB(n2215), .Q(\r[30][9] )
         );
  DFFARX1 \r_reg[30][8]  ( .D(n1016), .CLK(clk), .RSTB(n2215), .Q(\r[30][8] )
         );
  DFFARX1 \r_reg[30][7]  ( .D(n1015), .CLK(clk), .RSTB(n2215), .Q(\r[30][7] )
         );
  DFFARX1 \r_reg[30][6]  ( .D(n1014), .CLK(clk), .RSTB(n2215), .Q(\r[30][6] )
         );
  DFFARX1 \r_reg[30][5]  ( .D(n1013), .CLK(clk), .RSTB(n2215), .Q(\r[30][5] )
         );
  DFFARX1 \r_reg[30][4]  ( .D(n1012), .CLK(clk), .RSTB(n2215), .Q(\r[30][4] )
         );
  DFFARX1 \r_reg[30][3]  ( .D(n1011), .CLK(clk), .RSTB(n2216), .Q(\r[30][3] )
         );
  DFFARX1 \r_reg[30][2]  ( .D(n1010), .CLK(clk), .RSTB(n2216), .Q(\r[30][2] )
         );
  DFFARX1 \r_reg[30][1]  ( .D(n1009), .CLK(clk), .RSTB(n2216), .Q(\r[30][1] )
         );
  DFFARX1 \r_reg[30][0]  ( .D(n1008), .CLK(clk), .RSTB(n2216), .Q(\r[30][0] )
         );
  DFFARX1 \r_reg[29][31]  ( .D(n1007), .CLK(clk), .RSTB(n2216), .Q(\r[29][31] ) );
  DFFARX1 \r_reg[29][30]  ( .D(n1006), .CLK(clk), .RSTB(n2216), .Q(\r[29][30] ) );
  DFFARX1 \r_reg[29][29]  ( .D(n1005), .CLK(clk), .RSTB(n2216), .Q(\r[29][29] ) );
  DFFARX1 \r_reg[29][28]  ( .D(n1004), .CLK(clk), .RSTB(n2216), .Q(\r[29][28] ) );
  DFFARX1 \r_reg[29][27]  ( .D(n1003), .CLK(clk), .RSTB(n2216), .Q(\r[29][27] ) );
  DFFARX1 \r_reg[29][26]  ( .D(n1002), .CLK(clk), .RSTB(n2216), .Q(\r[29][26] ) );
  DFFARX1 \r_reg[29][25]  ( .D(n1001), .CLK(clk), .RSTB(n2216), .Q(\r[29][25] ) );
  DFFARX1 \r_reg[29][24]  ( .D(n1000), .CLK(clk), .RSTB(n2216), .Q(\r[29][24] ) );
  DFFARX1 \r_reg[29][23]  ( .D(n999), .CLK(clk), .RSTB(n2217), .Q(\r[29][23] )
         );
  DFFARX1 \r_reg[29][22]  ( .D(n998), .CLK(clk), .RSTB(n2217), .Q(\r[29][22] )
         );
  DFFARX1 \r_reg[29][21]  ( .D(n997), .CLK(clk), .RSTB(n2217), .Q(\r[29][21] )
         );
  DFFARX1 \r_reg[29][20]  ( .D(n996), .CLK(clk), .RSTB(n2217), .Q(\r[29][20] )
         );
  DFFARX1 \r_reg[29][19]  ( .D(n995), .CLK(clk), .RSTB(n2217), .Q(\r[29][19] )
         );
  DFFARX1 \r_reg[29][18]  ( .D(n994), .CLK(clk), .RSTB(n2217), .Q(\r[29][18] )
         );
  DFFARX1 \r_reg[29][17]  ( .D(n993), .CLK(clk), .RSTB(n2217), .Q(\r[29][17] )
         );
  DFFARX1 \r_reg[29][16]  ( .D(n992), .CLK(clk), .RSTB(n2217), .Q(\r[29][16] )
         );
  DFFARX1 \r_reg[29][15]  ( .D(n991), .CLK(clk), .RSTB(n2217), .Q(\r[29][15] )
         );
  DFFARX1 \r_reg[29][14]  ( .D(n990), .CLK(clk), .RSTB(n2217), .Q(\r[29][14] )
         );
  DFFARX1 \r_reg[29][13]  ( .D(n989), .CLK(clk), .RSTB(n2217), .Q(\r[29][13] )
         );
  DFFARX1 \r_reg[29][12]  ( .D(n988), .CLK(clk), .RSTB(n2217), .Q(\r[29][12] )
         );
  DFFARX1 \r_reg[29][11]  ( .D(n987), .CLK(clk), .RSTB(n2218), .Q(\r[29][11] )
         );
  DFFARX1 \r_reg[29][10]  ( .D(n986), .CLK(clk), .RSTB(n2218), .Q(\r[29][10] )
         );
  DFFARX1 \r_reg[29][9]  ( .D(n985), .CLK(clk), .RSTB(n2218), .Q(\r[29][9] )
         );
  DFFARX1 \r_reg[29][8]  ( .D(n984), .CLK(clk), .RSTB(n2218), .Q(\r[29][8] )
         );
  DFFARX1 \r_reg[29][7]  ( .D(n983), .CLK(clk), .RSTB(n2218), .Q(\r[29][7] )
         );
  DFFARX1 \r_reg[29][6]  ( .D(n982), .CLK(clk), .RSTB(n2218), .Q(\r[29][6] )
         );
  DFFARX1 \r_reg[29][5]  ( .D(n981), .CLK(clk), .RSTB(n2218), .Q(\r[29][5] )
         );
  DFFARX1 \r_reg[29][4]  ( .D(n980), .CLK(clk), .RSTB(n2218), .Q(\r[29][4] )
         );
  DFFARX1 \r_reg[29][3]  ( .D(n979), .CLK(clk), .RSTB(n2218), .Q(\r[29][3] )
         );
  DFFARX1 \r_reg[29][2]  ( .D(n978), .CLK(clk), .RSTB(n2218), .Q(\r[29][2] )
         );
  DFFARX1 \r_reg[29][1]  ( .D(n977), .CLK(clk), .RSTB(n2218), .Q(\r[29][1] )
         );
  DFFARX1 \r_reg[29][0]  ( .D(n976), .CLK(clk), .RSTB(n2218), .Q(\r[29][0] )
         );
  DFFARX1 \r_reg[28][31]  ( .D(n975), .CLK(clk), .RSTB(n2219), .Q(\r[28][31] )
         );
  DFFARX1 \r_reg[28][30]  ( .D(n974), .CLK(clk), .RSTB(n2219), .Q(\r[28][30] )
         );
  DFFARX1 \r_reg[28][29]  ( .D(n973), .CLK(clk), .RSTB(n2219), .Q(\r[28][29] )
         );
  DFFARX1 \r_reg[28][28]  ( .D(n972), .CLK(clk), .RSTB(n2219), .Q(\r[28][28] )
         );
  DFFARX1 \r_reg[28][27]  ( .D(n971), .CLK(clk), .RSTB(n2219), .Q(\r[28][27] )
         );
  DFFARX1 \r_reg[28][26]  ( .D(n970), .CLK(clk), .RSTB(n2219), .Q(\r[28][26] )
         );
  DFFARX1 \r_reg[28][25]  ( .D(n969), .CLK(clk), .RSTB(n2219), .Q(\r[28][25] )
         );
  DFFARX1 \r_reg[28][24]  ( .D(n968), .CLK(clk), .RSTB(n2219), .Q(\r[28][24] )
         );
  DFFARX1 \r_reg[28][23]  ( .D(n967), .CLK(clk), .RSTB(n2219), .Q(\r[28][23] )
         );
  DFFARX1 \r_reg[28][22]  ( .D(n966), .CLK(clk), .RSTB(n2219), .Q(\r[28][22] )
         );
  DFFARX1 \r_reg[28][21]  ( .D(n965), .CLK(clk), .RSTB(n2219), .Q(\r[28][21] )
         );
  DFFARX1 \r_reg[28][20]  ( .D(n964), .CLK(clk), .RSTB(n2219), .Q(\r[28][20] )
         );
  DFFARX1 \r_reg[28][19]  ( .D(n963), .CLK(clk), .RSTB(n2220), .Q(\r[28][19] )
         );
  DFFARX1 \r_reg[28][18]  ( .D(n962), .CLK(clk), .RSTB(n2220), .Q(\r[28][18] )
         );
  DFFARX1 \r_reg[28][17]  ( .D(n961), .CLK(clk), .RSTB(n2220), .Q(\r[28][17] )
         );
  DFFARX1 \r_reg[28][16]  ( .D(n960), .CLK(clk), .RSTB(n2220), .Q(\r[28][16] )
         );
  DFFARX1 \r_reg[28][15]  ( .D(n959), .CLK(clk), .RSTB(n2220), .Q(\r[28][15] )
         );
  DFFARX1 \r_reg[28][14]  ( .D(n958), .CLK(clk), .RSTB(n2220), .Q(\r[28][14] )
         );
  DFFARX1 \r_reg[28][13]  ( .D(n957), .CLK(clk), .RSTB(n2220), .Q(\r[28][13] )
         );
  DFFARX1 \r_reg[28][12]  ( .D(n956), .CLK(clk), .RSTB(n2220), .Q(\r[28][12] )
         );
  DFFARX1 \r_reg[28][11]  ( .D(n955), .CLK(clk), .RSTB(n2220), .Q(\r[28][11] )
         );
  DFFARX1 \r_reg[28][10]  ( .D(n954), .CLK(clk), .RSTB(n2220), .Q(\r[28][10] )
         );
  DFFARX1 \r_reg[28][9]  ( .D(n953), .CLK(clk), .RSTB(n2220), .Q(\r[28][9] )
         );
  DFFARX1 \r_reg[28][8]  ( .D(n952), .CLK(clk), .RSTB(n2220), .Q(\r[28][8] )
         );
  DFFARX1 \r_reg[28][7]  ( .D(n951), .CLK(clk), .RSTB(n2221), .Q(\r[28][7] )
         );
  DFFARX1 \r_reg[28][6]  ( .D(n950), .CLK(clk), .RSTB(n2221), .Q(\r[28][6] )
         );
  DFFARX1 \r_reg[28][5]  ( .D(n949), .CLK(clk), .RSTB(n2221), .Q(\r[28][5] )
         );
  DFFARX1 \r_reg[28][4]  ( .D(n948), .CLK(clk), .RSTB(n2221), .Q(\r[28][4] )
         );
  DFFARX1 \r_reg[28][3]  ( .D(n947), .CLK(clk), .RSTB(n2221), .Q(\r[28][3] )
         );
  DFFARX1 \r_reg[28][2]  ( .D(n946), .CLK(clk), .RSTB(n2221), .Q(\r[28][2] )
         );
  DFFARX1 \r_reg[28][1]  ( .D(n945), .CLK(clk), .RSTB(n2221), .Q(\r[28][1] )
         );
  DFFARX1 \r_reg[28][0]  ( .D(n944), .CLK(clk), .RSTB(n2221), .Q(\r[28][0] )
         );
  DFFARX1 \r_reg[27][31]  ( .D(n943), .CLK(clk), .RSTB(n2221), .Q(\r[27][31] )
         );
  DFFARX1 \r_reg[27][30]  ( .D(n942), .CLK(clk), .RSTB(n2221), .Q(\r[27][30] )
         );
  DFFARX1 \r_reg[27][29]  ( .D(n941), .CLK(clk), .RSTB(n2221), .Q(\r[27][29] )
         );
  DFFARX1 \r_reg[27][28]  ( .D(n940), .CLK(clk), .RSTB(n2221), .Q(\r[27][28] )
         );
  DFFARX1 \r_reg[27][27]  ( .D(n939), .CLK(clk), .RSTB(n2222), .Q(\r[27][27] )
         );
  DFFARX1 \r_reg[27][26]  ( .D(n938), .CLK(clk), .RSTB(n2222), .Q(\r[27][26] )
         );
  DFFARX1 \r_reg[27][25]  ( .D(n937), .CLK(clk), .RSTB(n2222), .Q(\r[27][25] )
         );
  DFFARX1 \r_reg[27][24]  ( .D(n936), .CLK(clk), .RSTB(n2222), .Q(\r[27][24] )
         );
  DFFARX1 \r_reg[27][23]  ( .D(n935), .CLK(clk), .RSTB(n2222), .Q(\r[27][23] )
         );
  DFFARX1 \r_reg[27][22]  ( .D(n934), .CLK(clk), .RSTB(n2222), .Q(\r[27][22] )
         );
  DFFARX1 \r_reg[27][21]  ( .D(n933), .CLK(clk), .RSTB(n2222), .Q(\r[27][21] )
         );
  DFFARX1 \r_reg[27][20]  ( .D(n932), .CLK(clk), .RSTB(n2222), .Q(\r[27][20] )
         );
  DFFARX1 \r_reg[27][19]  ( .D(n931), .CLK(clk), .RSTB(n2222), .Q(\r[27][19] )
         );
  DFFARX1 \r_reg[27][18]  ( .D(n930), .CLK(clk), .RSTB(n2222), .Q(\r[27][18] )
         );
  DFFARX1 \r_reg[27][17]  ( .D(n929), .CLK(clk), .RSTB(n2222), .Q(\r[27][17] )
         );
  DFFARX1 \r_reg[27][16]  ( .D(n928), .CLK(clk), .RSTB(n2222), .Q(\r[27][16] )
         );
  DFFARX1 \r_reg[27][15]  ( .D(n927), .CLK(clk), .RSTB(n2223), .Q(\r[27][15] )
         );
  DFFARX1 \r_reg[27][14]  ( .D(n926), .CLK(clk), .RSTB(n2223), .Q(\r[27][14] )
         );
  DFFARX1 \r_reg[27][13]  ( .D(n925), .CLK(clk), .RSTB(n2223), .Q(\r[27][13] )
         );
  DFFARX1 \r_reg[27][12]  ( .D(n924), .CLK(clk), .RSTB(n2223), .Q(\r[27][12] )
         );
  DFFARX1 \r_reg[27][11]  ( .D(n923), .CLK(clk), .RSTB(n2223), .Q(\r[27][11] )
         );
  DFFARX1 \r_reg[27][10]  ( .D(n922), .CLK(clk), .RSTB(n2223), .Q(\r[27][10] )
         );
  DFFARX1 \r_reg[27][9]  ( .D(n921), .CLK(clk), .RSTB(n2223), .Q(\r[27][9] )
         );
  DFFARX1 \r_reg[27][8]  ( .D(n920), .CLK(clk), .RSTB(n2223), .Q(\r[27][8] )
         );
  DFFARX1 \r_reg[27][7]  ( .D(n919), .CLK(clk), .RSTB(n2223), .Q(\r[27][7] )
         );
  DFFARX1 \r_reg[27][6]  ( .D(n918), .CLK(clk), .RSTB(n2223), .Q(\r[27][6] )
         );
  DFFARX1 \r_reg[27][5]  ( .D(n917), .CLK(clk), .RSTB(n2223), .Q(\r[27][5] )
         );
  DFFARX1 \r_reg[27][4]  ( .D(n916), .CLK(clk), .RSTB(n2223), .Q(\r[27][4] )
         );
  DFFARX1 \r_reg[27][3]  ( .D(n915), .CLK(clk), .RSTB(n2224), .Q(\r[27][3] )
         );
  DFFARX1 \r_reg[27][2]  ( .D(n914), .CLK(clk), .RSTB(n2224), .Q(\r[27][2] )
         );
  DFFARX1 \r_reg[27][1]  ( .D(n913), .CLK(clk), .RSTB(n2224), .Q(\r[27][1] )
         );
  DFFARX1 \r_reg[27][0]  ( .D(n912), .CLK(clk), .RSTB(n2224), .Q(\r[27][0] )
         );
  DFFARX1 \r_reg[26][31]  ( .D(n911), .CLK(clk), .RSTB(n2224), .Q(\r[26][31] )
         );
  DFFARX1 \r_reg[26][30]  ( .D(n910), .CLK(clk), .RSTB(n2224), .Q(\r[26][30] )
         );
  DFFARX1 \r_reg[26][29]  ( .D(n909), .CLK(clk), .RSTB(n2224), .Q(\r[26][29] )
         );
  DFFARX1 \r_reg[26][28]  ( .D(n908), .CLK(clk), .RSTB(n2224), .Q(\r[26][28] )
         );
  DFFARX1 \r_reg[26][27]  ( .D(n907), .CLK(clk), .RSTB(n2224), .Q(\r[26][27] )
         );
  DFFARX1 \r_reg[26][26]  ( .D(n906), .CLK(clk), .RSTB(n2224), .Q(\r[26][26] )
         );
  DFFARX1 \r_reg[26][25]  ( .D(n905), .CLK(clk), .RSTB(n2224), .Q(\r[26][25] )
         );
  DFFARX1 \r_reg[26][24]  ( .D(n904), .CLK(clk), .RSTB(n2224), .Q(\r[26][24] )
         );
  DFFARX1 \r_reg[26][23]  ( .D(n903), .CLK(clk), .RSTB(n2225), .Q(\r[26][23] )
         );
  DFFARX1 \r_reg[26][22]  ( .D(n902), .CLK(clk), .RSTB(n2225), .Q(\r[26][22] )
         );
  DFFARX1 \r_reg[26][21]  ( .D(n901), .CLK(clk), .RSTB(n2225), .Q(\r[26][21] )
         );
  DFFARX1 \r_reg[26][20]  ( .D(n900), .CLK(clk), .RSTB(n2225), .Q(\r[26][20] )
         );
  DFFARX1 \r_reg[26][19]  ( .D(n899), .CLK(clk), .RSTB(n2225), .Q(\r[26][19] )
         );
  DFFARX1 \r_reg[26][18]  ( .D(n898), .CLK(clk), .RSTB(n2225), .Q(\r[26][18] )
         );
  DFFARX1 \r_reg[26][17]  ( .D(n897), .CLK(clk), .RSTB(n2225), .Q(\r[26][17] )
         );
  DFFARX1 \r_reg[26][16]  ( .D(n896), .CLK(clk), .RSTB(n2225), .Q(\r[26][16] )
         );
  DFFARX1 \r_reg[26][15]  ( .D(n895), .CLK(clk), .RSTB(n2225), .Q(\r[26][15] )
         );
  DFFARX1 \r_reg[26][14]  ( .D(n894), .CLK(clk), .RSTB(n2225), .Q(\r[26][14] )
         );
  DFFARX1 \r_reg[26][13]  ( .D(n893), .CLK(clk), .RSTB(n2225), .Q(\r[26][13] )
         );
  DFFARX1 \r_reg[26][12]  ( .D(n892), .CLK(clk), .RSTB(n2225), .Q(\r[26][12] )
         );
  DFFARX1 \r_reg[26][11]  ( .D(n891), .CLK(clk), .RSTB(n2226), .Q(\r[26][11] )
         );
  DFFARX1 \r_reg[26][10]  ( .D(n890), .CLK(clk), .RSTB(n2226), .Q(\r[26][10] )
         );
  DFFARX1 \r_reg[26][9]  ( .D(n889), .CLK(clk), .RSTB(n2226), .Q(\r[26][9] )
         );
  DFFARX1 \r_reg[26][8]  ( .D(n888), .CLK(clk), .RSTB(n2226), .Q(\r[26][8] )
         );
  DFFARX1 \r_reg[26][7]  ( .D(n887), .CLK(clk), .RSTB(n2226), .Q(\r[26][7] )
         );
  DFFARX1 \r_reg[26][6]  ( .D(n886), .CLK(clk), .RSTB(n2226), .Q(\r[26][6] )
         );
  DFFARX1 \r_reg[26][5]  ( .D(n885), .CLK(clk), .RSTB(n2226), .Q(\r[26][5] )
         );
  DFFARX1 \r_reg[26][4]  ( .D(n884), .CLK(clk), .RSTB(n2226), .Q(\r[26][4] )
         );
  DFFARX1 \r_reg[26][3]  ( .D(n883), .CLK(clk), .RSTB(n2226), .Q(\r[26][3] )
         );
  DFFARX1 \r_reg[26][2]  ( .D(n882), .CLK(clk), .RSTB(n2226), .Q(\r[26][2] )
         );
  DFFARX1 \r_reg[26][1]  ( .D(n881), .CLK(clk), .RSTB(n2226), .Q(\r[26][1] )
         );
  DFFARX1 \r_reg[26][0]  ( .D(n880), .CLK(clk), .RSTB(n2226), .Q(\r[26][0] )
         );
  DFFARX1 \r_reg[25][31]  ( .D(n879), .CLK(clk), .RSTB(n2227), .Q(\r[25][31] )
         );
  DFFARX1 \r_reg[25][30]  ( .D(n878), .CLK(clk), .RSTB(n2227), .Q(\r[25][30] )
         );
  DFFARX1 \r_reg[25][29]  ( .D(n877), .CLK(clk), .RSTB(n2227), .Q(\r[25][29] )
         );
  DFFARX1 \r_reg[25][28]  ( .D(n876), .CLK(clk), .RSTB(n2227), .Q(\r[25][28] )
         );
  DFFARX1 \r_reg[25][27]  ( .D(n875), .CLK(clk), .RSTB(n2227), .Q(\r[25][27] )
         );
  DFFARX1 \r_reg[25][26]  ( .D(n874), .CLK(clk), .RSTB(n2227), .Q(\r[25][26] )
         );
  DFFARX1 \r_reg[25][25]  ( .D(n873), .CLK(clk), .RSTB(n2227), .Q(\r[25][25] )
         );
  DFFARX1 \r_reg[25][24]  ( .D(n872), .CLK(clk), .RSTB(n2227), .Q(\r[25][24] )
         );
  DFFARX1 \r_reg[25][23]  ( .D(n871), .CLK(clk), .RSTB(n2227), .Q(\r[25][23] )
         );
  DFFARX1 \r_reg[25][22]  ( .D(n870), .CLK(clk), .RSTB(n2227), .Q(\r[25][22] )
         );
  DFFARX1 \r_reg[25][21]  ( .D(n869), .CLK(clk), .RSTB(n2227), .Q(\r[25][21] )
         );
  DFFARX1 \r_reg[25][20]  ( .D(n868), .CLK(clk), .RSTB(n2227), .Q(\r[25][20] )
         );
  DFFARX1 \r_reg[25][19]  ( .D(n867), .CLK(clk), .RSTB(n2228), .Q(\r[25][19] )
         );
  DFFARX1 \r_reg[25][18]  ( .D(n866), .CLK(clk), .RSTB(n2228), .Q(\r[25][18] )
         );
  DFFARX1 \r_reg[25][17]  ( .D(n865), .CLK(clk), .RSTB(n2228), .Q(\r[25][17] )
         );
  DFFARX1 \r_reg[25][16]  ( .D(n864), .CLK(clk), .RSTB(n2228), .Q(\r[25][16] )
         );
  DFFARX1 \r_reg[25][15]  ( .D(n863), .CLK(clk), .RSTB(n2228), .Q(\r[25][15] )
         );
  DFFARX1 \r_reg[25][14]  ( .D(n862), .CLK(clk), .RSTB(n2228), .Q(\r[25][14] )
         );
  DFFARX1 \r_reg[25][13]  ( .D(n861), .CLK(clk), .RSTB(n2228), .Q(\r[25][13] )
         );
  DFFARX1 \r_reg[25][12]  ( .D(n860), .CLK(clk), .RSTB(n2228), .Q(\r[25][12] )
         );
  DFFARX1 \r_reg[25][11]  ( .D(n859), .CLK(clk), .RSTB(n2228), .Q(\r[25][11] )
         );
  DFFARX1 \r_reg[25][10]  ( .D(n858), .CLK(clk), .RSTB(n2228), .Q(\r[25][10] )
         );
  DFFARX1 \r_reg[25][9]  ( .D(n857), .CLK(clk), .RSTB(n2228), .Q(\r[25][9] )
         );
  DFFARX1 \r_reg[25][8]  ( .D(n856), .CLK(clk), .RSTB(n2228), .Q(\r[25][8] )
         );
  DFFARX1 \r_reg[25][7]  ( .D(n855), .CLK(clk), .RSTB(n2229), .Q(\r[25][7] )
         );
  DFFARX1 \r_reg[25][6]  ( .D(n854), .CLK(clk), .RSTB(n2229), .Q(\r[25][6] )
         );
  DFFARX1 \r_reg[25][5]  ( .D(n853), .CLK(clk), .RSTB(n2229), .Q(\r[25][5] )
         );
  DFFARX1 \r_reg[25][4]  ( .D(n852), .CLK(clk), .RSTB(n2229), .Q(\r[25][4] )
         );
  DFFARX1 \r_reg[25][3]  ( .D(n851), .CLK(clk), .RSTB(n2229), .Q(\r[25][3] )
         );
  DFFARX1 \r_reg[25][2]  ( .D(n850), .CLK(clk), .RSTB(n2229), .Q(\r[25][2] )
         );
  DFFARX1 \r_reg[25][1]  ( .D(n849), .CLK(clk), .RSTB(n2229), .Q(\r[25][1] )
         );
  DFFARX1 \r_reg[25][0]  ( .D(n848), .CLK(clk), .RSTB(n2229), .Q(\r[25][0] )
         );
  DFFARX1 \r_reg[24][31]  ( .D(n847), .CLK(clk), .RSTB(n2229), .Q(\r[24][31] )
         );
  DFFARX1 \r_reg[24][30]  ( .D(n846), .CLK(clk), .RSTB(n2229), .Q(\r[24][30] )
         );
  DFFARX1 \r_reg[24][29]  ( .D(n845), .CLK(clk), .RSTB(n2229), .Q(\r[24][29] )
         );
  DFFARX1 \r_reg[24][28]  ( .D(n844), .CLK(clk), .RSTB(n2229), .Q(\r[24][28] )
         );
  DFFARX1 \r_reg[24][27]  ( .D(n843), .CLK(clk), .RSTB(n2230), .Q(\r[24][27] )
         );
  DFFARX1 \r_reg[24][26]  ( .D(n842), .CLK(clk), .RSTB(n2230), .Q(\r[24][26] )
         );
  DFFARX1 \r_reg[24][25]  ( .D(n841), .CLK(clk), .RSTB(n2230), .Q(\r[24][25] )
         );
  DFFARX1 \r_reg[24][24]  ( .D(n840), .CLK(clk), .RSTB(n2230), .Q(\r[24][24] )
         );
  DFFARX1 \r_reg[24][23]  ( .D(n839), .CLK(clk), .RSTB(n2230), .Q(\r[24][23] )
         );
  DFFARX1 \r_reg[24][22]  ( .D(n838), .CLK(clk), .RSTB(n2230), .Q(\r[24][22] )
         );
  DFFARX1 \r_reg[24][21]  ( .D(n837), .CLK(clk), .RSTB(n2230), .Q(\r[24][21] )
         );
  DFFARX1 \r_reg[24][20]  ( .D(n836), .CLK(clk), .RSTB(n2230), .Q(\r[24][20] )
         );
  DFFARX1 \r_reg[24][19]  ( .D(n835), .CLK(clk), .RSTB(n2230), .Q(\r[24][19] )
         );
  DFFARX1 \r_reg[24][18]  ( .D(n834), .CLK(clk), .RSTB(n2230), .Q(\r[24][18] )
         );
  DFFARX1 \r_reg[24][17]  ( .D(n833), .CLK(clk), .RSTB(n2230), .Q(\r[24][17] )
         );
  DFFARX1 \r_reg[24][16]  ( .D(n832), .CLK(clk), .RSTB(n2230), .Q(\r[24][16] )
         );
  DFFARX1 \r_reg[24][15]  ( .D(n831), .CLK(clk), .RSTB(n2231), .Q(\r[24][15] )
         );
  DFFARX1 \r_reg[24][14]  ( .D(n830), .CLK(clk), .RSTB(n2231), .Q(\r[24][14] )
         );
  DFFARX1 \r_reg[24][13]  ( .D(n829), .CLK(clk), .RSTB(n2231), .Q(\r[24][13] )
         );
  DFFARX1 \r_reg[24][12]  ( .D(n828), .CLK(clk), .RSTB(n2231), .Q(\r[24][12] )
         );
  DFFARX1 \r_reg[24][11]  ( .D(n827), .CLK(clk), .RSTB(n2231), .Q(\r[24][11] )
         );
  DFFARX1 \r_reg[24][10]  ( .D(n826), .CLK(clk), .RSTB(n2231), .Q(\r[24][10] )
         );
  DFFARX1 \r_reg[24][9]  ( .D(n825), .CLK(clk), .RSTB(n2231), .Q(\r[24][9] )
         );
  DFFARX1 \r_reg[24][8]  ( .D(n824), .CLK(clk), .RSTB(n2231), .Q(\r[24][8] )
         );
  DFFARX1 \r_reg[24][7]  ( .D(n823), .CLK(clk), .RSTB(n2231), .Q(\r[24][7] )
         );
  DFFARX1 \r_reg[24][6]  ( .D(n822), .CLK(clk), .RSTB(n2231), .Q(\r[24][6] )
         );
  DFFARX1 \r_reg[24][5]  ( .D(n821), .CLK(clk), .RSTB(n2231), .Q(\r[24][5] )
         );
  DFFARX1 \r_reg[24][4]  ( .D(n820), .CLK(clk), .RSTB(n2231), .Q(\r[24][4] )
         );
  DFFARX1 \r_reg[24][3]  ( .D(n819), .CLK(clk), .RSTB(n2232), .Q(\r[24][3] )
         );
  DFFARX1 \r_reg[24][2]  ( .D(n818), .CLK(clk), .RSTB(n2232), .Q(\r[24][2] )
         );
  DFFARX1 \r_reg[24][1]  ( .D(n817), .CLK(clk), .RSTB(n2232), .Q(\r[24][1] )
         );
  DFFARX1 \r_reg[24][0]  ( .D(n816), .CLK(clk), .RSTB(n2232), .Q(\r[24][0] )
         );
  DFFARX1 \r_reg[23][31]  ( .D(n815), .CLK(clk), .RSTB(n2232), .Q(\r[23][31] )
         );
  DFFARX1 \r_reg[23][30]  ( .D(n814), .CLK(clk), .RSTB(n2232), .Q(\r[23][30] )
         );
  DFFARX1 \r_reg[23][29]  ( .D(n813), .CLK(clk), .RSTB(n2232), .Q(\r[23][29] )
         );
  DFFARX1 \r_reg[23][28]  ( .D(n812), .CLK(clk), .RSTB(n2232), .Q(\r[23][28] )
         );
  DFFARX1 \r_reg[23][27]  ( .D(n811), .CLK(clk), .RSTB(n2232), .Q(\r[23][27] )
         );
  DFFARX1 \r_reg[23][26]  ( .D(n810), .CLK(clk), .RSTB(n2232), .Q(\r[23][26] )
         );
  DFFARX1 \r_reg[23][25]  ( .D(n809), .CLK(clk), .RSTB(n2232), .Q(\r[23][25] )
         );
  DFFARX1 \r_reg[23][24]  ( .D(n808), .CLK(clk), .RSTB(n2232), .Q(\r[23][24] )
         );
  DFFARX1 \r_reg[23][23]  ( .D(n807), .CLK(clk), .RSTB(n2233), .Q(\r[23][23] )
         );
  DFFARX1 \r_reg[23][22]  ( .D(n806), .CLK(clk), .RSTB(n2233), .Q(\r[23][22] )
         );
  DFFARX1 \r_reg[23][21]  ( .D(n805), .CLK(clk), .RSTB(n2233), .Q(\r[23][21] )
         );
  DFFARX1 \r_reg[23][20]  ( .D(n804), .CLK(clk), .RSTB(n2233), .Q(\r[23][20] )
         );
  DFFARX1 \r_reg[23][19]  ( .D(n803), .CLK(clk), .RSTB(n2233), .Q(\r[23][19] )
         );
  DFFARX1 \r_reg[23][18]  ( .D(n802), .CLK(clk), .RSTB(n2233), .Q(\r[23][18] )
         );
  DFFARX1 \r_reg[23][17]  ( .D(n801), .CLK(clk), .RSTB(n2233), .Q(\r[23][17] )
         );
  DFFARX1 \r_reg[23][16]  ( .D(n800), .CLK(clk), .RSTB(n2233), .Q(\r[23][16] )
         );
  DFFARX1 \r_reg[23][15]  ( .D(n799), .CLK(clk), .RSTB(n2233), .Q(\r[23][15] )
         );
  DFFARX1 \r_reg[23][14]  ( .D(n798), .CLK(clk), .RSTB(n2233), .Q(\r[23][14] )
         );
  DFFARX1 \r_reg[23][13]  ( .D(n797), .CLK(clk), .RSTB(n2233), .Q(\r[23][13] )
         );
  DFFARX1 \r_reg[23][12]  ( .D(n796), .CLK(clk), .RSTB(n2233), .Q(\r[23][12] )
         );
  DFFARX1 \r_reg[23][11]  ( .D(n795), .CLK(clk), .RSTB(n2234), .Q(\r[23][11] )
         );
  DFFARX1 \r_reg[23][10]  ( .D(n794), .CLK(clk), .RSTB(n2234), .Q(\r[23][10] )
         );
  DFFARX1 \r_reg[23][9]  ( .D(n793), .CLK(clk), .RSTB(n2234), .Q(\r[23][9] )
         );
  DFFARX1 \r_reg[23][8]  ( .D(n792), .CLK(clk), .RSTB(n2234), .Q(\r[23][8] )
         );
  DFFARX1 \r_reg[23][7]  ( .D(n791), .CLK(clk), .RSTB(n2234), .Q(\r[23][7] )
         );
  DFFARX1 \r_reg[23][6]  ( .D(n790), .CLK(clk), .RSTB(n2234), .Q(\r[23][6] )
         );
  DFFARX1 \r_reg[23][5]  ( .D(n789), .CLK(clk), .RSTB(n2234), .Q(\r[23][5] )
         );
  DFFARX1 \r_reg[23][4]  ( .D(n788), .CLK(clk), .RSTB(n2234), .Q(\r[23][4] )
         );
  DFFARX1 \r_reg[23][3]  ( .D(n787), .CLK(clk), .RSTB(n2234), .Q(\r[23][3] )
         );
  DFFARX1 \r_reg[23][2]  ( .D(n786), .CLK(clk), .RSTB(n2234), .Q(\r[23][2] )
         );
  DFFARX1 \r_reg[23][1]  ( .D(n785), .CLK(clk), .RSTB(n2234), .Q(\r[23][1] )
         );
  DFFARX1 \r_reg[23][0]  ( .D(n784), .CLK(clk), .RSTB(n2234), .Q(\r[23][0] )
         );
  DFFARX1 \r_reg[22][31]  ( .D(n783), .CLK(clk), .RSTB(n2235), .Q(\r[22][31] )
         );
  DFFARX1 \r_reg[22][30]  ( .D(n782), .CLK(clk), .RSTB(n2235), .Q(\r[22][30] )
         );
  DFFARX1 \r_reg[22][29]  ( .D(n781), .CLK(clk), .RSTB(n2235), .Q(\r[22][29] )
         );
  DFFARX1 \r_reg[22][28]  ( .D(n780), .CLK(clk), .RSTB(n2235), .Q(\r[22][28] )
         );
  DFFARX1 \r_reg[22][27]  ( .D(n779), .CLK(clk), .RSTB(n2235), .Q(\r[22][27] )
         );
  DFFARX1 \r_reg[22][26]  ( .D(n778), .CLK(clk), .RSTB(n2235), .Q(\r[22][26] )
         );
  DFFARX1 \r_reg[22][25]  ( .D(n777), .CLK(clk), .RSTB(n2235), .Q(\r[22][25] )
         );
  DFFARX1 \r_reg[22][24]  ( .D(n776), .CLK(clk), .RSTB(n2235), .Q(\r[22][24] )
         );
  DFFARX1 \r_reg[22][23]  ( .D(n775), .CLK(clk), .RSTB(n2235), .Q(\r[22][23] )
         );
  DFFARX1 \r_reg[22][22]  ( .D(n774), .CLK(clk), .RSTB(n2235), .Q(\r[22][22] )
         );
  DFFARX1 \r_reg[22][21]  ( .D(n773), .CLK(clk), .RSTB(n2235), .Q(\r[22][21] )
         );
  DFFARX1 \r_reg[22][20]  ( .D(n772), .CLK(clk), .RSTB(n2235), .Q(\r[22][20] )
         );
  DFFARX1 \r_reg[22][19]  ( .D(n771), .CLK(clk), .RSTB(n2236), .Q(\r[22][19] )
         );
  DFFARX1 \r_reg[22][18]  ( .D(n770), .CLK(clk), .RSTB(n2236), .Q(\r[22][18] )
         );
  DFFARX1 \r_reg[22][17]  ( .D(n769), .CLK(clk), .RSTB(n2236), .Q(\r[22][17] )
         );
  DFFARX1 \r_reg[22][16]  ( .D(n768), .CLK(clk), .RSTB(n2236), .Q(\r[22][16] )
         );
  DFFARX1 \r_reg[22][15]  ( .D(n767), .CLK(clk), .RSTB(n2236), .Q(\r[22][15] )
         );
  DFFARX1 \r_reg[22][14]  ( .D(n766), .CLK(clk), .RSTB(n2236), .Q(\r[22][14] )
         );
  DFFARX1 \r_reg[22][13]  ( .D(n765), .CLK(clk), .RSTB(n2236), .Q(\r[22][13] )
         );
  DFFARX1 \r_reg[22][12]  ( .D(n764), .CLK(clk), .RSTB(n2236), .Q(\r[22][12] )
         );
  DFFARX1 \r_reg[22][11]  ( .D(n763), .CLK(clk), .RSTB(n2236), .Q(\r[22][11] )
         );
  DFFARX1 \r_reg[22][10]  ( .D(n762), .CLK(clk), .RSTB(n2236), .Q(\r[22][10] )
         );
  DFFARX1 \r_reg[22][9]  ( .D(n761), .CLK(clk), .RSTB(n2236), .Q(\r[22][9] )
         );
  DFFARX1 \r_reg[22][8]  ( .D(n760), .CLK(clk), .RSTB(n2236), .Q(\r[22][8] )
         );
  DFFARX1 \r_reg[22][7]  ( .D(n759), .CLK(clk), .RSTB(n2237), .Q(\r[22][7] )
         );
  DFFARX1 \r_reg[22][6]  ( .D(n758), .CLK(clk), .RSTB(n2237), .Q(\r[22][6] )
         );
  DFFARX1 \r_reg[22][5]  ( .D(n757), .CLK(clk), .RSTB(n2237), .Q(\r[22][5] )
         );
  DFFARX1 \r_reg[22][4]  ( .D(n756), .CLK(clk), .RSTB(n2237), .Q(\r[22][4] )
         );
  DFFARX1 \r_reg[22][3]  ( .D(n755), .CLK(clk), .RSTB(n2237), .Q(\r[22][3] )
         );
  DFFARX1 \r_reg[22][2]  ( .D(n754), .CLK(clk), .RSTB(n2237), .Q(\r[22][2] )
         );
  DFFARX1 \r_reg[22][1]  ( .D(n753), .CLK(clk), .RSTB(n2237), .Q(\r[22][1] )
         );
  DFFARX1 \r_reg[22][0]  ( .D(n752), .CLK(clk), .RSTB(n2237), .Q(\r[22][0] )
         );
  DFFARX1 \r_reg[21][31]  ( .D(n751), .CLK(clk), .RSTB(n2237), .Q(\r[21][31] )
         );
  DFFARX1 \r_reg[21][30]  ( .D(n750), .CLK(clk), .RSTB(n2237), .Q(\r[21][30] )
         );
  DFFARX1 \r_reg[21][29]  ( .D(n749), .CLK(clk), .RSTB(n2237), .Q(\r[21][29] )
         );
  DFFARX1 \r_reg[21][28]  ( .D(n748), .CLK(clk), .RSTB(n2237), .Q(\r[21][28] )
         );
  DFFARX1 \r_reg[21][27]  ( .D(n747), .CLK(clk), .RSTB(n2238), .Q(\r[21][27] )
         );
  DFFARX1 \r_reg[21][26]  ( .D(n746), .CLK(clk), .RSTB(n2238), .Q(\r[21][26] )
         );
  DFFARX1 \r_reg[21][25]  ( .D(n745), .CLK(clk), .RSTB(n2238), .Q(\r[21][25] )
         );
  DFFARX1 \r_reg[21][24]  ( .D(n744), .CLK(clk), .RSTB(n2238), .Q(\r[21][24] )
         );
  DFFARX1 \r_reg[21][23]  ( .D(n743), .CLK(clk), .RSTB(n2238), .Q(\r[21][23] )
         );
  DFFARX1 \r_reg[21][22]  ( .D(n742), .CLK(clk), .RSTB(n2238), .Q(\r[21][22] )
         );
  DFFARX1 \r_reg[21][21]  ( .D(n741), .CLK(clk), .RSTB(n2238), .Q(\r[21][21] )
         );
  DFFARX1 \r_reg[21][20]  ( .D(n740), .CLK(clk), .RSTB(n2238), .Q(\r[21][20] )
         );
  DFFARX1 \r_reg[21][19]  ( .D(n739), .CLK(clk), .RSTB(n2238), .Q(\r[21][19] )
         );
  DFFARX1 \r_reg[21][18]  ( .D(n738), .CLK(clk), .RSTB(n2238), .Q(\r[21][18] )
         );
  DFFARX1 \r_reg[21][17]  ( .D(n737), .CLK(clk), .RSTB(n2238), .Q(\r[21][17] )
         );
  DFFARX1 \r_reg[21][16]  ( .D(n736), .CLK(clk), .RSTB(n2238), .Q(\r[21][16] )
         );
  DFFARX1 \r_reg[21][15]  ( .D(n735), .CLK(clk), .RSTB(n2239), .Q(\r[21][15] )
         );
  DFFARX1 \r_reg[21][14]  ( .D(n734), .CLK(clk), .RSTB(n2239), .Q(\r[21][14] )
         );
  DFFARX1 \r_reg[21][13]  ( .D(n733), .CLK(clk), .RSTB(n2239), .Q(\r[21][13] )
         );
  DFFARX1 \r_reg[21][12]  ( .D(n732), .CLK(clk), .RSTB(n2239), .Q(\r[21][12] )
         );
  DFFARX1 \r_reg[21][11]  ( .D(n731), .CLK(clk), .RSTB(n2239), .Q(\r[21][11] )
         );
  DFFARX1 \r_reg[21][10]  ( .D(n730), .CLK(clk), .RSTB(n2239), .Q(\r[21][10] )
         );
  DFFARX1 \r_reg[21][9]  ( .D(n729), .CLK(clk), .RSTB(n2239), .Q(\r[21][9] )
         );
  DFFARX1 \r_reg[21][8]  ( .D(n728), .CLK(clk), .RSTB(n2239), .Q(\r[21][8] )
         );
  DFFARX1 \r_reg[21][7]  ( .D(n727), .CLK(clk), .RSTB(n2239), .Q(\r[21][7] )
         );
  DFFARX1 \r_reg[21][6]  ( .D(n726), .CLK(clk), .RSTB(n2239), .Q(\r[21][6] )
         );
  DFFARX1 \r_reg[21][5]  ( .D(n725), .CLK(clk), .RSTB(n2239), .Q(\r[21][5] )
         );
  DFFARX1 \r_reg[21][4]  ( .D(n724), .CLK(clk), .RSTB(n2239), .Q(\r[21][4] )
         );
  DFFARX1 \r_reg[21][3]  ( .D(n723), .CLK(clk), .RSTB(n2240), .Q(\r[21][3] )
         );
  DFFARX1 \r_reg[21][2]  ( .D(n722), .CLK(clk), .RSTB(n2240), .Q(\r[21][2] )
         );
  DFFARX1 \r_reg[21][1]  ( .D(n721), .CLK(clk), .RSTB(n2240), .Q(\r[21][1] )
         );
  DFFARX1 \r_reg[21][0]  ( .D(n720), .CLK(clk), .RSTB(n2240), .Q(\r[21][0] )
         );
  DFFARX1 \r_reg[20][31]  ( .D(n719), .CLK(clk), .RSTB(n2240), .Q(\r[20][31] )
         );
  DFFARX1 \r_reg[20][30]  ( .D(n718), .CLK(clk), .RSTB(n2240), .Q(\r[20][30] )
         );
  DFFARX1 \r_reg[20][29]  ( .D(n717), .CLK(clk), .RSTB(n2240), .Q(\r[20][29] )
         );
  DFFARX1 \r_reg[20][28]  ( .D(n716), .CLK(clk), .RSTB(n2240), .Q(\r[20][28] )
         );
  DFFARX1 \r_reg[20][27]  ( .D(n715), .CLK(clk), .RSTB(n2240), .Q(\r[20][27] )
         );
  DFFARX1 \r_reg[20][26]  ( .D(n714), .CLK(clk), .RSTB(n2240), .Q(\r[20][26] )
         );
  DFFARX1 \r_reg[20][25]  ( .D(n713), .CLK(clk), .RSTB(n2240), .Q(\r[20][25] )
         );
  DFFARX1 \r_reg[20][24]  ( .D(n712), .CLK(clk), .RSTB(n2240), .Q(\r[20][24] )
         );
  DFFARX1 \r_reg[20][23]  ( .D(n711), .CLK(clk), .RSTB(n2241), .Q(\r[20][23] )
         );
  DFFARX1 \r_reg[20][22]  ( .D(n710), .CLK(clk), .RSTB(n2241), .Q(\r[20][22] )
         );
  DFFARX1 \r_reg[20][21]  ( .D(n709), .CLK(clk), .RSTB(n2241), .Q(\r[20][21] )
         );
  DFFARX1 \r_reg[20][20]  ( .D(n708), .CLK(clk), .RSTB(n2241), .Q(\r[20][20] )
         );
  DFFARX1 \r_reg[20][19]  ( .D(n707), .CLK(clk), .RSTB(n2241), .Q(\r[20][19] )
         );
  DFFARX1 \r_reg[20][18]  ( .D(n706), .CLK(clk), .RSTB(n2241), .Q(\r[20][18] )
         );
  DFFARX1 \r_reg[20][17]  ( .D(n705), .CLK(clk), .RSTB(n2241), .Q(\r[20][17] )
         );
  DFFARX1 \r_reg[20][16]  ( .D(n704), .CLK(clk), .RSTB(n2241), .Q(\r[20][16] )
         );
  DFFARX1 \r_reg[20][15]  ( .D(n703), .CLK(clk), .RSTB(n2241), .Q(\r[20][15] )
         );
  DFFARX1 \r_reg[20][14]  ( .D(n702), .CLK(clk), .RSTB(n2241), .Q(\r[20][14] )
         );
  DFFARX1 \r_reg[20][13]  ( .D(n701), .CLK(clk), .RSTB(n2241), .Q(\r[20][13] )
         );
  DFFARX1 \r_reg[20][12]  ( .D(n700), .CLK(clk), .RSTB(n2241), .Q(\r[20][12] )
         );
  DFFARX1 \r_reg[20][11]  ( .D(n699), .CLK(clk), .RSTB(n2242), .Q(\r[20][11] )
         );
  DFFARX1 \r_reg[20][10]  ( .D(n698), .CLK(clk), .RSTB(n2242), .Q(\r[20][10] )
         );
  DFFARX1 \r_reg[20][9]  ( .D(n697), .CLK(clk), .RSTB(n2242), .Q(\r[20][9] )
         );
  DFFARX1 \r_reg[20][8]  ( .D(n696), .CLK(clk), .RSTB(n2242), .Q(\r[20][8] )
         );
  DFFARX1 \r_reg[20][7]  ( .D(n695), .CLK(clk), .RSTB(n2242), .Q(\r[20][7] )
         );
  DFFARX1 \r_reg[20][6]  ( .D(n694), .CLK(clk), .RSTB(n2242), .Q(\r[20][6] )
         );
  DFFARX1 \r_reg[20][5]  ( .D(n693), .CLK(clk), .RSTB(n2242), .Q(\r[20][5] )
         );
  DFFARX1 \r_reg[20][4]  ( .D(n692), .CLK(clk), .RSTB(n2242), .Q(\r[20][4] )
         );
  DFFARX1 \r_reg[20][3]  ( .D(n691), .CLK(clk), .RSTB(n2242), .Q(\r[20][3] )
         );
  DFFARX1 \r_reg[20][2]  ( .D(n690), .CLK(clk), .RSTB(n2242), .Q(\r[20][2] )
         );
  DFFARX1 \r_reg[20][1]  ( .D(n689), .CLK(clk), .RSTB(n2242), .Q(\r[20][1] )
         );
  DFFARX1 \r_reg[20][0]  ( .D(n688), .CLK(clk), .RSTB(n2242), .Q(\r[20][0] )
         );
  DFFARX1 \r_reg[19][31]  ( .D(n687), .CLK(clk), .RSTB(n2243), .Q(\r[19][31] )
         );
  DFFARX1 \r_reg[19][30]  ( .D(n686), .CLK(clk), .RSTB(n2243), .Q(\r[19][30] )
         );
  DFFARX1 \r_reg[19][29]  ( .D(n685), .CLK(clk), .RSTB(n2243), .Q(\r[19][29] )
         );
  DFFARX1 \r_reg[19][28]  ( .D(n684), .CLK(clk), .RSTB(n2243), .Q(\r[19][28] )
         );
  DFFARX1 \r_reg[19][27]  ( .D(n683), .CLK(clk), .RSTB(n2243), .Q(\r[19][27] )
         );
  DFFARX1 \r_reg[19][26]  ( .D(n682), .CLK(clk), .RSTB(n2243), .Q(\r[19][26] )
         );
  DFFARX1 \r_reg[19][25]  ( .D(n681), .CLK(clk), .RSTB(n2243), .Q(\r[19][25] )
         );
  DFFARX1 \r_reg[19][24]  ( .D(n680), .CLK(clk), .RSTB(n2243), .Q(\r[19][24] )
         );
  DFFARX1 \r_reg[19][23]  ( .D(n679), .CLK(clk), .RSTB(n2243), .Q(\r[19][23] )
         );
  DFFARX1 \r_reg[19][22]  ( .D(n678), .CLK(clk), .RSTB(n2243), .Q(\r[19][22] )
         );
  DFFARX1 \r_reg[19][21]  ( .D(n677), .CLK(clk), .RSTB(n2243), .Q(\r[19][21] )
         );
  DFFARX1 \r_reg[19][20]  ( .D(n676), .CLK(clk), .RSTB(n2243), .Q(\r[19][20] )
         );
  DFFARX1 \r_reg[19][19]  ( .D(n675), .CLK(clk), .RSTB(n2244), .Q(\r[19][19] )
         );
  DFFARX1 \r_reg[19][18]  ( .D(n674), .CLK(clk), .RSTB(n2244), .Q(\r[19][18] )
         );
  DFFARX1 \r_reg[19][17]  ( .D(n673), .CLK(clk), .RSTB(n2244), .Q(\r[19][17] )
         );
  DFFARX1 \r_reg[19][16]  ( .D(n672), .CLK(clk), .RSTB(n2244), .Q(\r[19][16] )
         );
  DFFARX1 \r_reg[19][15]  ( .D(n671), .CLK(clk), .RSTB(n2244), .Q(\r[19][15] )
         );
  DFFARX1 \r_reg[19][14]  ( .D(n670), .CLK(clk), .RSTB(n2244), .Q(\r[19][14] )
         );
  DFFARX1 \r_reg[19][13]  ( .D(n669), .CLK(clk), .RSTB(n2244), .Q(\r[19][13] )
         );
  DFFARX1 \r_reg[19][12]  ( .D(n668), .CLK(clk), .RSTB(n2244), .Q(\r[19][12] )
         );
  DFFARX1 \r_reg[19][11]  ( .D(n667), .CLK(clk), .RSTB(n2244), .Q(\r[19][11] )
         );
  DFFARX1 \r_reg[19][10]  ( .D(n666), .CLK(clk), .RSTB(n2244), .Q(\r[19][10] )
         );
  DFFARX1 \r_reg[19][9]  ( .D(n665), .CLK(clk), .RSTB(n2244), .Q(\r[19][9] )
         );
  DFFARX1 \r_reg[19][8]  ( .D(n664), .CLK(clk), .RSTB(n2244), .Q(\r[19][8] )
         );
  DFFARX1 \r_reg[19][7]  ( .D(n663), .CLK(clk), .RSTB(n2245), .Q(\r[19][7] )
         );
  DFFARX1 \r_reg[19][6]  ( .D(n662), .CLK(clk), .RSTB(n2245), .Q(\r[19][6] )
         );
  DFFARX1 \r_reg[19][5]  ( .D(n661), .CLK(clk), .RSTB(n2245), .Q(\r[19][5] )
         );
  DFFARX1 \r_reg[19][4]  ( .D(n660), .CLK(clk), .RSTB(n2245), .Q(\r[19][4] )
         );
  DFFARX1 \r_reg[19][3]  ( .D(n659), .CLK(clk), .RSTB(n2245), .Q(\r[19][3] )
         );
  DFFARX1 \r_reg[19][2]  ( .D(n658), .CLK(clk), .RSTB(n2245), .Q(\r[19][2] )
         );
  DFFARX1 \r_reg[19][1]  ( .D(n657), .CLK(clk), .RSTB(n2245), .Q(\r[19][1] )
         );
  DFFARX1 \r_reg[19][0]  ( .D(n656), .CLK(clk), .RSTB(n2245), .Q(\r[19][0] )
         );
  DFFARX1 \r_reg[18][31]  ( .D(n655), .CLK(clk), .RSTB(n2245), .Q(\r[18][31] )
         );
  DFFARX1 \r_reg[18][30]  ( .D(n654), .CLK(clk), .RSTB(n2245), .Q(\r[18][30] )
         );
  DFFARX1 \r_reg[18][29]  ( .D(n653), .CLK(clk), .RSTB(n2245), .Q(\r[18][29] )
         );
  DFFARX1 \r_reg[18][28]  ( .D(n652), .CLK(clk), .RSTB(n2245), .Q(\r[18][28] )
         );
  DFFARX1 \r_reg[18][27]  ( .D(n651), .CLK(clk), .RSTB(n2246), .Q(\r[18][27] )
         );
  DFFARX1 \r_reg[18][26]  ( .D(n650), .CLK(clk), .RSTB(n2246), .Q(\r[18][26] )
         );
  DFFARX1 \r_reg[18][25]  ( .D(n649), .CLK(clk), .RSTB(n2246), .Q(\r[18][25] )
         );
  DFFARX1 \r_reg[18][24]  ( .D(n648), .CLK(clk), .RSTB(n2246), .Q(\r[18][24] )
         );
  DFFARX1 \r_reg[18][23]  ( .D(n647), .CLK(clk), .RSTB(n2246), .Q(\r[18][23] )
         );
  DFFARX1 \r_reg[18][22]  ( .D(n646), .CLK(clk), .RSTB(n2246), .Q(\r[18][22] )
         );
  DFFARX1 \r_reg[18][21]  ( .D(n645), .CLK(clk), .RSTB(n2246), .Q(\r[18][21] )
         );
  DFFARX1 \r_reg[18][20]  ( .D(n644), .CLK(clk), .RSTB(n2246), .Q(\r[18][20] )
         );
  DFFARX1 \r_reg[18][19]  ( .D(n643), .CLK(clk), .RSTB(n2246), .Q(\r[18][19] )
         );
  DFFARX1 \r_reg[18][18]  ( .D(n642), .CLK(clk), .RSTB(n2246), .Q(\r[18][18] )
         );
  DFFARX1 \r_reg[18][17]  ( .D(n641), .CLK(clk), .RSTB(n2246), .Q(\r[18][17] )
         );
  DFFARX1 \r_reg[18][16]  ( .D(n640), .CLK(clk), .RSTB(n2246), .Q(\r[18][16] )
         );
  DFFARX1 \r_reg[18][15]  ( .D(n639), .CLK(clk), .RSTB(n2247), .Q(\r[18][15] )
         );
  DFFARX1 \r_reg[18][14]  ( .D(n638), .CLK(clk), .RSTB(n2247), .Q(\r[18][14] )
         );
  DFFARX1 \r_reg[18][13]  ( .D(n637), .CLK(clk), .RSTB(n2247), .Q(\r[18][13] )
         );
  DFFARX1 \r_reg[18][12]  ( .D(n636), .CLK(clk), .RSTB(n2247), .Q(\r[18][12] )
         );
  DFFARX1 \r_reg[18][11]  ( .D(n635), .CLK(clk), .RSTB(n2247), .Q(\r[18][11] )
         );
  DFFARX1 \r_reg[18][10]  ( .D(n634), .CLK(clk), .RSTB(n2247), .Q(\r[18][10] )
         );
  DFFARX1 \r_reg[18][9]  ( .D(n633), .CLK(clk), .RSTB(n2247), .Q(\r[18][9] )
         );
  DFFARX1 \r_reg[18][8]  ( .D(n632), .CLK(clk), .RSTB(n2247), .Q(\r[18][8] )
         );
  DFFARX1 \r_reg[18][7]  ( .D(n631), .CLK(clk), .RSTB(n2247), .Q(\r[18][7] )
         );
  DFFARX1 \r_reg[18][6]  ( .D(n630), .CLK(clk), .RSTB(n2247), .Q(\r[18][6] )
         );
  DFFARX1 \r_reg[18][5]  ( .D(n629), .CLK(clk), .RSTB(n2247), .Q(\r[18][5] )
         );
  DFFARX1 \r_reg[18][4]  ( .D(n628), .CLK(clk), .RSTB(n2247), .Q(\r[18][4] )
         );
  DFFARX1 \r_reg[18][3]  ( .D(n627), .CLK(clk), .RSTB(n2248), .Q(\r[18][3] )
         );
  DFFARX1 \r_reg[18][2]  ( .D(n626), .CLK(clk), .RSTB(n2248), .Q(\r[18][2] )
         );
  DFFARX1 \r_reg[18][1]  ( .D(n625), .CLK(clk), .RSTB(n2248), .Q(\r[18][1] )
         );
  DFFARX1 \r_reg[18][0]  ( .D(n624), .CLK(clk), .RSTB(n2248), .Q(\r[18][0] )
         );
  DFFARX1 \r_reg[17][31]  ( .D(n623), .CLK(clk), .RSTB(n2248), .Q(\r[17][31] )
         );
  DFFARX1 \r_reg[17][30]  ( .D(n622), .CLK(clk), .RSTB(n2248), .Q(\r[17][30] )
         );
  DFFARX1 \r_reg[17][29]  ( .D(n621), .CLK(clk), .RSTB(n2248), .Q(\r[17][29] )
         );
  DFFARX1 \r_reg[17][28]  ( .D(n620), .CLK(clk), .RSTB(n2248), .Q(\r[17][28] )
         );
  DFFARX1 \r_reg[17][27]  ( .D(n619), .CLK(clk), .RSTB(n2248), .Q(\r[17][27] )
         );
  DFFARX1 \r_reg[17][26]  ( .D(n618), .CLK(clk), .RSTB(n2248), .Q(\r[17][26] )
         );
  DFFARX1 \r_reg[17][25]  ( .D(n617), .CLK(clk), .RSTB(n2248), .Q(\r[17][25] )
         );
  DFFARX1 \r_reg[17][24]  ( .D(n616), .CLK(clk), .RSTB(n2248), .Q(\r[17][24] )
         );
  DFFARX1 \r_reg[17][23]  ( .D(n615), .CLK(clk), .RSTB(n2249), .Q(\r[17][23] )
         );
  DFFARX1 \r_reg[17][22]  ( .D(n614), .CLK(clk), .RSTB(n2249), .Q(\r[17][22] )
         );
  DFFARX1 \r_reg[17][21]  ( .D(n613), .CLK(clk), .RSTB(n2249), .Q(\r[17][21] )
         );
  DFFARX1 \r_reg[17][20]  ( .D(n612), .CLK(clk), .RSTB(n2249), .Q(\r[17][20] )
         );
  DFFARX1 \r_reg[17][19]  ( .D(n611), .CLK(clk), .RSTB(n2249), .Q(\r[17][19] )
         );
  DFFARX1 \r_reg[17][18]  ( .D(n610), .CLK(clk), .RSTB(n2249), .Q(\r[17][18] )
         );
  DFFARX1 \r_reg[17][17]  ( .D(n609), .CLK(clk), .RSTB(n2249), .Q(\r[17][17] )
         );
  DFFARX1 \r_reg[17][16]  ( .D(n608), .CLK(clk), .RSTB(n2249), .Q(\r[17][16] )
         );
  DFFARX1 \r_reg[17][15]  ( .D(n607), .CLK(clk), .RSTB(n2249), .Q(\r[17][15] )
         );
  DFFARX1 \r_reg[17][14]  ( .D(n606), .CLK(clk), .RSTB(n2249), .Q(\r[17][14] )
         );
  DFFARX1 \r_reg[17][13]  ( .D(n605), .CLK(clk), .RSTB(n2249), .Q(\r[17][13] )
         );
  DFFARX1 \r_reg[17][12]  ( .D(n604), .CLK(clk), .RSTB(n2249), .Q(\r[17][12] )
         );
  DFFARX1 \r_reg[17][11]  ( .D(n603), .CLK(clk), .RSTB(n2250), .Q(\r[17][11] )
         );
  DFFARX1 \r_reg[17][10]  ( .D(n602), .CLK(clk), .RSTB(n2250), .Q(\r[17][10] )
         );
  DFFARX1 \r_reg[17][9]  ( .D(n601), .CLK(clk), .RSTB(n2250), .Q(\r[17][9] )
         );
  DFFARX1 \r_reg[17][8]  ( .D(n600), .CLK(clk), .RSTB(n2250), .Q(\r[17][8] )
         );
  DFFARX1 \r_reg[17][7]  ( .D(n599), .CLK(clk), .RSTB(n2250), .Q(\r[17][7] )
         );
  DFFARX1 \r_reg[17][6]  ( .D(n598), .CLK(clk), .RSTB(n2250), .Q(\r[17][6] )
         );
  DFFARX1 \r_reg[17][5]  ( .D(n597), .CLK(clk), .RSTB(n2250), .Q(\r[17][5] )
         );
  DFFARX1 \r_reg[17][4]  ( .D(n596), .CLK(clk), .RSTB(n2250), .Q(\r[17][4] )
         );
  DFFARX1 \r_reg[17][3]  ( .D(n595), .CLK(clk), .RSTB(n2250), .Q(\r[17][3] )
         );
  DFFARX1 \r_reg[17][2]  ( .D(n594), .CLK(clk), .RSTB(n2250), .Q(\r[17][2] )
         );
  DFFARX1 \r_reg[17][1]  ( .D(n593), .CLK(clk), .RSTB(n2250), .Q(\r[17][1] )
         );
  DFFARX1 \r_reg[17][0]  ( .D(n592), .CLK(clk), .RSTB(n2250), .Q(\r[17][0] )
         );
  DFFARX1 \r_reg[16][31]  ( .D(n591), .CLK(clk), .RSTB(n2251), .Q(\r[16][31] )
         );
  DFFARX1 \r_reg[16][30]  ( .D(n590), .CLK(clk), .RSTB(n2251), .Q(\r[16][30] )
         );
  DFFARX1 \r_reg[16][29]  ( .D(n589), .CLK(clk), .RSTB(n2251), .Q(\r[16][29] )
         );
  DFFARX1 \r_reg[16][28]  ( .D(n588), .CLK(clk), .RSTB(n2251), .Q(\r[16][28] )
         );
  DFFARX1 \r_reg[16][27]  ( .D(n587), .CLK(clk), .RSTB(n2251), .Q(\r[16][27] )
         );
  DFFARX1 \r_reg[16][26]  ( .D(n586), .CLK(clk), .RSTB(n2251), .Q(\r[16][26] )
         );
  DFFARX1 \r_reg[16][25]  ( .D(n585), .CLK(clk), .RSTB(n2251), .Q(\r[16][25] )
         );
  DFFARX1 \r_reg[16][24]  ( .D(n584), .CLK(clk), .RSTB(n2251), .Q(\r[16][24] )
         );
  DFFARX1 \r_reg[16][23]  ( .D(n583), .CLK(clk), .RSTB(n2251), .Q(\r[16][23] )
         );
  DFFARX1 \r_reg[16][22]  ( .D(n582), .CLK(clk), .RSTB(n2251), .Q(\r[16][22] )
         );
  DFFARX1 \r_reg[16][21]  ( .D(n581), .CLK(clk), .RSTB(n2251), .Q(\r[16][21] )
         );
  DFFARX1 \r_reg[16][20]  ( .D(n580), .CLK(clk), .RSTB(n2251), .Q(\r[16][20] )
         );
  DFFARX1 \r_reg[16][19]  ( .D(n579), .CLK(clk), .RSTB(n2252), .Q(\r[16][19] )
         );
  DFFARX1 \r_reg[16][18]  ( .D(n578), .CLK(clk), .RSTB(n2252), .Q(\r[16][18] )
         );
  DFFARX1 \r_reg[16][17]  ( .D(n577), .CLK(clk), .RSTB(n2252), .Q(\r[16][17] )
         );
  DFFARX1 \r_reg[16][16]  ( .D(n576), .CLK(clk), .RSTB(n2252), .Q(\r[16][16] )
         );
  DFFARX1 \r_reg[16][15]  ( .D(n575), .CLK(clk), .RSTB(n2252), .Q(\r[16][15] )
         );
  DFFARX1 \r_reg[16][14]  ( .D(n574), .CLK(clk), .RSTB(n2252), .Q(\r[16][14] )
         );
  DFFARX1 \r_reg[16][13]  ( .D(n573), .CLK(clk), .RSTB(n2252), .Q(\r[16][13] )
         );
  DFFARX1 \r_reg[16][12]  ( .D(n572), .CLK(clk), .RSTB(n2252), .Q(\r[16][12] )
         );
  DFFARX1 \r_reg[16][11]  ( .D(n571), .CLK(clk), .RSTB(n2252), .Q(\r[16][11] )
         );
  DFFARX1 \r_reg[16][10]  ( .D(n570), .CLK(clk), .RSTB(n2252), .Q(\r[16][10] )
         );
  DFFARX1 \r_reg[16][9]  ( .D(n569), .CLK(clk), .RSTB(n2252), .Q(\r[16][9] )
         );
  DFFARX1 \r_reg[16][8]  ( .D(n568), .CLK(clk), .RSTB(n2252), .Q(\r[16][8] )
         );
  DFFARX1 \r_reg[16][7]  ( .D(n567), .CLK(clk), .RSTB(n2253), .Q(\r[16][7] )
         );
  DFFARX1 \r_reg[16][6]  ( .D(n566), .CLK(clk), .RSTB(n2253), .Q(\r[16][6] )
         );
  DFFARX1 \r_reg[16][5]  ( .D(n565), .CLK(clk), .RSTB(n2253), .Q(\r[16][5] )
         );
  DFFARX1 \r_reg[16][4]  ( .D(n564), .CLK(clk), .RSTB(n2253), .Q(\r[16][4] )
         );
  DFFARX1 \r_reg[16][3]  ( .D(n563), .CLK(clk), .RSTB(n2253), .Q(\r[16][3] )
         );
  DFFARX1 \r_reg[16][2]  ( .D(n562), .CLK(clk), .RSTB(n2253), .Q(\r[16][2] )
         );
  DFFARX1 \r_reg[16][1]  ( .D(n561), .CLK(clk), .RSTB(n2253), .Q(\r[16][1] )
         );
  DFFARX1 \r_reg[16][0]  ( .D(n560), .CLK(clk), .RSTB(n2253), .Q(\r[16][0] )
         );
  DFFARX1 \r_reg[15][31]  ( .D(n559), .CLK(clk), .RSTB(n2253), .Q(\r[15][31] )
         );
  DFFARX1 \r_reg[15][30]  ( .D(n558), .CLK(clk), .RSTB(n2253), .Q(\r[15][30] )
         );
  DFFARX1 \r_reg[15][29]  ( .D(n557), .CLK(clk), .RSTB(n2253), .Q(\r[15][29] )
         );
  DFFARX1 \r_reg[15][28]  ( .D(n556), .CLK(clk), .RSTB(n2253), .Q(\r[15][28] )
         );
  DFFARX1 \r_reg[15][27]  ( .D(n555), .CLK(clk), .RSTB(n2254), .Q(\r[15][27] )
         );
  DFFARX1 \r_reg[15][26]  ( .D(n554), .CLK(clk), .RSTB(n2254), .Q(\r[15][26] )
         );
  DFFARX1 \r_reg[15][25]  ( .D(n553), .CLK(clk), .RSTB(n2254), .Q(\r[15][25] )
         );
  DFFARX1 \r_reg[15][24]  ( .D(n552), .CLK(clk), .RSTB(n2254), .Q(\r[15][24] )
         );
  DFFARX1 \r_reg[15][23]  ( .D(n551), .CLK(clk), .RSTB(n2254), .Q(\r[15][23] )
         );
  DFFARX1 \r_reg[15][22]  ( .D(n550), .CLK(clk), .RSTB(n2254), .Q(\r[15][22] )
         );
  DFFARX1 \r_reg[15][21]  ( .D(n549), .CLK(clk), .RSTB(n2254), .Q(\r[15][21] )
         );
  DFFARX1 \r_reg[15][20]  ( .D(n548), .CLK(clk), .RSTB(n2254), .Q(\r[15][20] )
         );
  DFFARX1 \r_reg[15][19]  ( .D(n547), .CLK(clk), .RSTB(n2254), .Q(\r[15][19] )
         );
  DFFARX1 \r_reg[15][18]  ( .D(n546), .CLK(clk), .RSTB(n2254), .Q(\r[15][18] )
         );
  DFFARX1 \r_reg[15][17]  ( .D(n545), .CLK(clk), .RSTB(n2254), .Q(\r[15][17] )
         );
  DFFARX1 \r_reg[15][16]  ( .D(n544), .CLK(clk), .RSTB(n2254), .Q(\r[15][16] )
         );
  DFFARX1 \r_reg[15][15]  ( .D(n543), .CLK(clk), .RSTB(n2255), .Q(\r[15][15] )
         );
  DFFARX1 \r_reg[15][14]  ( .D(n542), .CLK(clk), .RSTB(n2255), .Q(\r[15][14] )
         );
  DFFARX1 \r_reg[15][13]  ( .D(n541), .CLK(clk), .RSTB(n2255), .Q(\r[15][13] )
         );
  DFFARX1 \r_reg[15][12]  ( .D(n540), .CLK(clk), .RSTB(n2255), .Q(\r[15][12] )
         );
  DFFARX1 \r_reg[15][11]  ( .D(n539), .CLK(clk), .RSTB(n2255), .Q(\r[15][11] )
         );
  DFFARX1 \r_reg[15][10]  ( .D(n538), .CLK(clk), .RSTB(n2255), .Q(\r[15][10] )
         );
  DFFARX1 \r_reg[15][9]  ( .D(n537), .CLK(clk), .RSTB(n2255), .Q(\r[15][9] )
         );
  DFFARX1 \r_reg[15][8]  ( .D(n536), .CLK(clk), .RSTB(n2255), .Q(\r[15][8] )
         );
  DFFARX1 \r_reg[15][7]  ( .D(n535), .CLK(clk), .RSTB(n2255), .Q(\r[15][7] )
         );
  DFFARX1 \r_reg[15][6]  ( .D(n534), .CLK(clk), .RSTB(n2255), .Q(\r[15][6] )
         );
  DFFARX1 \r_reg[15][5]  ( .D(n533), .CLK(clk), .RSTB(n2255), .Q(\r[15][5] )
         );
  DFFARX1 \r_reg[15][4]  ( .D(n532), .CLK(clk), .RSTB(n2255), .Q(\r[15][4] )
         );
  DFFARX1 \r_reg[15][3]  ( .D(n531), .CLK(clk), .RSTB(n2256), .Q(\r[15][3] )
         );
  DFFARX1 \r_reg[15][2]  ( .D(n530), .CLK(clk), .RSTB(n2256), .Q(\r[15][2] )
         );
  DFFARX1 \r_reg[15][1]  ( .D(n529), .CLK(clk), .RSTB(n2256), .Q(\r[15][1] )
         );
  DFFARX1 \r_reg[15][0]  ( .D(n528), .CLK(clk), .RSTB(n2256), .Q(\r[15][0] )
         );
  DFFARX1 \r_reg[14][31]  ( .D(n527), .CLK(clk), .RSTB(n2256), .Q(\r[14][31] )
         );
  DFFARX1 \r_reg[14][30]  ( .D(n526), .CLK(clk), .RSTB(n2256), .Q(\r[14][30] )
         );
  DFFARX1 \r_reg[14][29]  ( .D(n525), .CLK(clk), .RSTB(n2256), .Q(\r[14][29] )
         );
  DFFARX1 \r_reg[14][28]  ( .D(n524), .CLK(clk), .RSTB(n2256), .Q(\r[14][28] )
         );
  DFFARX1 \r_reg[14][27]  ( .D(n523), .CLK(clk), .RSTB(n2256), .Q(\r[14][27] )
         );
  DFFARX1 \r_reg[14][26]  ( .D(n522), .CLK(clk), .RSTB(n2256), .Q(\r[14][26] )
         );
  DFFARX1 \r_reg[14][25]  ( .D(n521), .CLK(clk), .RSTB(n2256), .Q(\r[14][25] )
         );
  DFFARX1 \r_reg[14][24]  ( .D(n520), .CLK(clk), .RSTB(n2256), .Q(\r[14][24] )
         );
  DFFARX1 \r_reg[14][23]  ( .D(n519), .CLK(clk), .RSTB(n2257), .Q(\r[14][23] )
         );
  DFFARX1 \r_reg[14][22]  ( .D(n518), .CLK(clk), .RSTB(n2257), .Q(\r[14][22] )
         );
  DFFARX1 \r_reg[14][21]  ( .D(n517), .CLK(clk), .RSTB(n2257), .Q(\r[14][21] )
         );
  DFFARX1 \r_reg[14][20]  ( .D(n516), .CLK(clk), .RSTB(n2257), .Q(\r[14][20] )
         );
  DFFARX1 \r_reg[14][19]  ( .D(n515), .CLK(clk), .RSTB(n2257), .Q(\r[14][19] )
         );
  DFFARX1 \r_reg[14][18]  ( .D(n514), .CLK(clk), .RSTB(n2257), .Q(\r[14][18] )
         );
  DFFARX1 \r_reg[14][17]  ( .D(n513), .CLK(clk), .RSTB(n2257), .Q(\r[14][17] )
         );
  DFFARX1 \r_reg[14][16]  ( .D(n512), .CLK(clk), .RSTB(n2257), .Q(\r[14][16] )
         );
  DFFARX1 \r_reg[14][15]  ( .D(n511), .CLK(clk), .RSTB(n2257), .Q(\r[14][15] )
         );
  DFFARX1 \r_reg[14][14]  ( .D(n510), .CLK(clk), .RSTB(n2257), .Q(\r[14][14] )
         );
  DFFARX1 \r_reg[14][13]  ( .D(n509), .CLK(clk), .RSTB(n2257), .Q(\r[14][13] )
         );
  DFFARX1 \r_reg[14][12]  ( .D(n508), .CLK(clk), .RSTB(n2257), .Q(\r[14][12] )
         );
  DFFARX1 \r_reg[14][11]  ( .D(n507), .CLK(clk), .RSTB(n2258), .Q(\r[14][11] )
         );
  DFFARX1 \r_reg[14][10]  ( .D(n506), .CLK(clk), .RSTB(n2258), .Q(\r[14][10] )
         );
  DFFARX1 \r_reg[14][9]  ( .D(n505), .CLK(clk), .RSTB(n2258), .Q(\r[14][9] )
         );
  DFFARX1 \r_reg[14][8]  ( .D(n504), .CLK(clk), .RSTB(n2258), .Q(\r[14][8] )
         );
  DFFARX1 \r_reg[14][7]  ( .D(n503), .CLK(clk), .RSTB(n2258), .Q(\r[14][7] )
         );
  DFFARX1 \r_reg[14][6]  ( .D(n502), .CLK(clk), .RSTB(n2258), .Q(\r[14][6] )
         );
  DFFARX1 \r_reg[14][5]  ( .D(n501), .CLK(clk), .RSTB(n2258), .Q(\r[14][5] )
         );
  DFFARX1 \r_reg[14][4]  ( .D(n500), .CLK(clk), .RSTB(n2258), .Q(\r[14][4] )
         );
  DFFARX1 \r_reg[14][3]  ( .D(n499), .CLK(clk), .RSTB(n2258), .Q(\r[14][3] )
         );
  DFFARX1 \r_reg[14][2]  ( .D(n498), .CLK(clk), .RSTB(n2258), .Q(\r[14][2] )
         );
  DFFARX1 \r_reg[14][1]  ( .D(n497), .CLK(clk), .RSTB(n2258), .Q(\r[14][1] )
         );
  DFFARX1 \r_reg[14][0]  ( .D(n496), .CLK(clk), .RSTB(n2258), .Q(\r[14][0] )
         );
  DFFARX1 \r_reg[13][31]  ( .D(n495), .CLK(clk), .RSTB(n2259), .Q(\r[13][31] )
         );
  DFFARX1 \r_reg[13][30]  ( .D(n494), .CLK(clk), .RSTB(n2259), .Q(\r[13][30] )
         );
  DFFARX1 \r_reg[13][29]  ( .D(n493), .CLK(clk), .RSTB(n2259), .Q(\r[13][29] )
         );
  DFFARX1 \r_reg[13][28]  ( .D(n492), .CLK(clk), .RSTB(n2259), .Q(\r[13][28] )
         );
  DFFARX1 \r_reg[13][27]  ( .D(n491), .CLK(clk), .RSTB(n2259), .Q(\r[13][27] )
         );
  DFFARX1 \r_reg[13][26]  ( .D(n490), .CLK(clk), .RSTB(n2259), .Q(\r[13][26] )
         );
  DFFARX1 \r_reg[13][25]  ( .D(n489), .CLK(clk), .RSTB(n2259), .Q(\r[13][25] )
         );
  DFFARX1 \r_reg[13][24]  ( .D(n488), .CLK(clk), .RSTB(n2259), .Q(\r[13][24] )
         );
  DFFARX1 \r_reg[13][23]  ( .D(n487), .CLK(clk), .RSTB(n2259), .Q(\r[13][23] )
         );
  DFFARX1 \r_reg[13][22]  ( .D(n486), .CLK(clk), .RSTB(n2259), .Q(\r[13][22] )
         );
  DFFARX1 \r_reg[13][21]  ( .D(n485), .CLK(clk), .RSTB(n2259), .Q(\r[13][21] )
         );
  DFFARX1 \r_reg[13][20]  ( .D(n484), .CLK(clk), .RSTB(n2259), .Q(\r[13][20] )
         );
  DFFARX1 \r_reg[13][19]  ( .D(n483), .CLK(clk), .RSTB(n2260), .Q(\r[13][19] )
         );
  DFFARX1 \r_reg[13][18]  ( .D(n482), .CLK(clk), .RSTB(n2260), .Q(\r[13][18] )
         );
  DFFARX1 \r_reg[13][17]  ( .D(n481), .CLK(clk), .RSTB(n2260), .Q(\r[13][17] )
         );
  DFFARX1 \r_reg[13][16]  ( .D(n480), .CLK(clk), .RSTB(n2260), .Q(\r[13][16] )
         );
  DFFARX1 \r_reg[13][15]  ( .D(n479), .CLK(clk), .RSTB(n2260), .Q(\r[13][15] )
         );
  DFFARX1 \r_reg[13][14]  ( .D(n478), .CLK(clk), .RSTB(n2260), .Q(\r[13][14] )
         );
  DFFARX1 \r_reg[13][13]  ( .D(n477), .CLK(clk), .RSTB(n2260), .Q(\r[13][13] )
         );
  DFFARX1 \r_reg[13][12]  ( .D(n476), .CLK(clk), .RSTB(n2260), .Q(\r[13][12] )
         );
  DFFARX1 \r_reg[13][11]  ( .D(n475), .CLK(clk), .RSTB(n2260), .Q(\r[13][11] )
         );
  DFFARX1 \r_reg[13][10]  ( .D(n474), .CLK(clk), .RSTB(n2260), .Q(\r[13][10] )
         );
  DFFARX1 \r_reg[13][9]  ( .D(n473), .CLK(clk), .RSTB(n2260), .Q(\r[13][9] )
         );
  DFFARX1 \r_reg[13][8]  ( .D(n472), .CLK(clk), .RSTB(n2260), .Q(\r[13][8] )
         );
  DFFARX1 \r_reg[13][7]  ( .D(n471), .CLK(clk), .RSTB(n2261), .Q(\r[13][7] )
         );
  DFFARX1 \r_reg[13][6]  ( .D(n470), .CLK(clk), .RSTB(n2261), .Q(\r[13][6] )
         );
  DFFARX1 \r_reg[13][5]  ( .D(n469), .CLK(clk), .RSTB(n2261), .Q(\r[13][5] )
         );
  DFFARX1 \r_reg[13][4]  ( .D(n468), .CLK(clk), .RSTB(n2261), .Q(\r[13][4] )
         );
  DFFARX1 \r_reg[13][3]  ( .D(n467), .CLK(clk), .RSTB(n2261), .Q(\r[13][3] )
         );
  DFFARX1 \r_reg[13][2]  ( .D(n466), .CLK(clk), .RSTB(n2261), .Q(\r[13][2] )
         );
  DFFARX1 \r_reg[13][1]  ( .D(n465), .CLK(clk), .RSTB(n2261), .Q(\r[13][1] )
         );
  DFFARX1 \r_reg[13][0]  ( .D(n464), .CLK(clk), .RSTB(n2261), .Q(\r[13][0] )
         );
  DFFARX1 \r_reg[12][31]  ( .D(n463), .CLK(clk), .RSTB(n2261), .Q(\r[12][31] )
         );
  DFFARX1 \r_reg[12][30]  ( .D(n462), .CLK(clk), .RSTB(n2261), .Q(\r[12][30] )
         );
  DFFARX1 \r_reg[12][29]  ( .D(n461), .CLK(clk), .RSTB(n2261), .Q(\r[12][29] )
         );
  DFFARX1 \r_reg[12][28]  ( .D(n460), .CLK(clk), .RSTB(n2261), .Q(\r[12][28] )
         );
  DFFARX1 \r_reg[12][27]  ( .D(n459), .CLK(clk), .RSTB(n2262), .Q(\r[12][27] )
         );
  DFFARX1 \r_reg[12][26]  ( .D(n458), .CLK(clk), .RSTB(n2262), .Q(\r[12][26] )
         );
  DFFARX1 \r_reg[12][25]  ( .D(n457), .CLK(clk), .RSTB(n2262), .Q(\r[12][25] )
         );
  DFFARX1 \r_reg[12][24]  ( .D(n456), .CLK(clk), .RSTB(n2262), .Q(\r[12][24] )
         );
  DFFARX1 \r_reg[12][23]  ( .D(n455), .CLK(clk), .RSTB(n2262), .Q(\r[12][23] )
         );
  DFFARX1 \r_reg[12][22]  ( .D(n454), .CLK(clk), .RSTB(n2262), .Q(\r[12][22] )
         );
  DFFARX1 \r_reg[12][21]  ( .D(n453), .CLK(clk), .RSTB(n2262), .Q(\r[12][21] )
         );
  DFFARX1 \r_reg[12][20]  ( .D(n452), .CLK(clk), .RSTB(n2262), .Q(\r[12][20] )
         );
  DFFARX1 \r_reg[12][19]  ( .D(n451), .CLK(clk), .RSTB(n2262), .Q(\r[12][19] )
         );
  DFFARX1 \r_reg[12][18]  ( .D(n450), .CLK(clk), .RSTB(n2262), .Q(\r[12][18] )
         );
  DFFARX1 \r_reg[12][17]  ( .D(n449), .CLK(clk), .RSTB(n2262), .Q(\r[12][17] )
         );
  DFFARX1 \r_reg[12][16]  ( .D(n448), .CLK(clk), .RSTB(n2262), .Q(\r[12][16] )
         );
  DFFARX1 \r_reg[12][15]  ( .D(n447), .CLK(clk), .RSTB(n2263), .Q(\r[12][15] )
         );
  DFFARX1 \r_reg[12][14]  ( .D(n446), .CLK(clk), .RSTB(n2263), .Q(\r[12][14] )
         );
  DFFARX1 \r_reg[12][13]  ( .D(n445), .CLK(clk), .RSTB(n2263), .Q(\r[12][13] )
         );
  DFFARX1 \r_reg[12][12]  ( .D(n444), .CLK(clk), .RSTB(n2263), .Q(\r[12][12] )
         );
  DFFARX1 \r_reg[12][11]  ( .D(n443), .CLK(clk), .RSTB(n2263), .Q(\r[12][11] )
         );
  DFFARX1 \r_reg[12][10]  ( .D(n442), .CLK(clk), .RSTB(n2263), .Q(\r[12][10] )
         );
  DFFARX1 \r_reg[12][9]  ( .D(n441), .CLK(clk), .RSTB(n2263), .Q(\r[12][9] )
         );
  DFFARX1 \r_reg[12][8]  ( .D(n440), .CLK(clk), .RSTB(n2263), .Q(\r[12][8] )
         );
  DFFARX1 \r_reg[12][7]  ( .D(n439), .CLK(clk), .RSTB(n2263), .Q(\r[12][7] )
         );
  DFFARX1 \r_reg[12][6]  ( .D(n438), .CLK(clk), .RSTB(n2263), .Q(\r[12][6] )
         );
  DFFARX1 \r_reg[12][5]  ( .D(n437), .CLK(clk), .RSTB(n2263), .Q(\r[12][5] )
         );
  DFFARX1 \r_reg[12][4]  ( .D(n436), .CLK(clk), .RSTB(n2263), .Q(\r[12][4] )
         );
  DFFARX1 \r_reg[12][3]  ( .D(n435), .CLK(clk), .RSTB(n2264), .Q(\r[12][3] )
         );
  DFFARX1 \r_reg[12][2]  ( .D(n434), .CLK(clk), .RSTB(n2264), .Q(\r[12][2] )
         );
  DFFARX1 \r_reg[12][1]  ( .D(n433), .CLK(clk), .RSTB(n2264), .Q(\r[12][1] )
         );
  DFFARX1 \r_reg[12][0]  ( .D(n432), .CLK(clk), .RSTB(n2264), .Q(\r[12][0] )
         );
  DFFARX1 \r_reg[11][31]  ( .D(n431), .CLK(clk), .RSTB(n2264), .Q(\r[11][31] )
         );
  DFFARX1 \r_reg[11][30]  ( .D(n430), .CLK(clk), .RSTB(n2264), .Q(\r[11][30] )
         );
  DFFARX1 \r_reg[11][29]  ( .D(n429), .CLK(clk), .RSTB(n2264), .Q(\r[11][29] )
         );
  DFFARX1 \r_reg[11][28]  ( .D(n428), .CLK(clk), .RSTB(n2264), .Q(\r[11][28] )
         );
  DFFARX1 \r_reg[11][27]  ( .D(n427), .CLK(clk), .RSTB(n2264), .Q(\r[11][27] )
         );
  DFFARX1 \r_reg[11][26]  ( .D(n426), .CLK(clk), .RSTB(n2264), .Q(\r[11][26] )
         );
  DFFARX1 \r_reg[11][25]  ( .D(n425), .CLK(clk), .RSTB(n2264), .Q(\r[11][25] )
         );
  DFFARX1 \r_reg[11][24]  ( .D(n424), .CLK(clk), .RSTB(n2264), .Q(\r[11][24] )
         );
  DFFARX1 \r_reg[11][23]  ( .D(n423), .CLK(clk), .RSTB(n2265), .Q(\r[11][23] )
         );
  DFFARX1 \r_reg[11][22]  ( .D(n422), .CLK(clk), .RSTB(n2265), .Q(\r[11][22] )
         );
  DFFARX1 \r_reg[11][21]  ( .D(n421), .CLK(clk), .RSTB(n2265), .Q(\r[11][21] )
         );
  DFFARX1 \r_reg[11][20]  ( .D(n420), .CLK(clk), .RSTB(n2265), .Q(\r[11][20] )
         );
  DFFARX1 \r_reg[11][19]  ( .D(n419), .CLK(clk), .RSTB(n2265), .Q(\r[11][19] )
         );
  DFFARX1 \r_reg[11][18]  ( .D(n418), .CLK(clk), .RSTB(n2265), .Q(\r[11][18] )
         );
  DFFARX1 \r_reg[11][17]  ( .D(n417), .CLK(clk), .RSTB(n2265), .Q(\r[11][17] )
         );
  DFFARX1 \r_reg[11][16]  ( .D(n416), .CLK(clk), .RSTB(n2265), .Q(\r[11][16] )
         );
  DFFARX1 \r_reg[11][15]  ( .D(n415), .CLK(clk), .RSTB(n2265), .Q(\r[11][15] )
         );
  DFFARX1 \r_reg[11][14]  ( .D(n414), .CLK(clk), .RSTB(n2265), .Q(\r[11][14] )
         );
  DFFARX1 \r_reg[11][13]  ( .D(n413), .CLK(clk), .RSTB(n2265), .Q(\r[11][13] )
         );
  DFFARX1 \r_reg[11][12]  ( .D(n412), .CLK(clk), .RSTB(n2265), .Q(\r[11][12] )
         );
  DFFARX1 \r_reg[11][11]  ( .D(n411), .CLK(clk), .RSTB(n2266), .Q(\r[11][11] )
         );
  DFFARX1 \r_reg[11][10]  ( .D(n410), .CLK(clk), .RSTB(n2266), .Q(\r[11][10] )
         );
  DFFARX1 \r_reg[11][9]  ( .D(n409), .CLK(clk), .RSTB(n2266), .Q(\r[11][9] )
         );
  DFFARX1 \r_reg[11][8]  ( .D(n408), .CLK(clk), .RSTB(n2266), .Q(\r[11][8] )
         );
  DFFARX1 \r_reg[11][7]  ( .D(n407), .CLK(clk), .RSTB(n2266), .Q(\r[11][7] )
         );
  DFFARX1 \r_reg[11][6]  ( .D(n406), .CLK(clk), .RSTB(n2266), .Q(\r[11][6] )
         );
  DFFARX1 \r_reg[11][5]  ( .D(n405), .CLK(clk), .RSTB(n2266), .Q(\r[11][5] )
         );
  DFFARX1 \r_reg[11][4]  ( .D(n404), .CLK(clk), .RSTB(n2266), .Q(\r[11][4] )
         );
  DFFARX1 \r_reg[11][3]  ( .D(n403), .CLK(clk), .RSTB(n2266), .Q(\r[11][3] )
         );
  DFFARX1 \r_reg[11][2]  ( .D(n402), .CLK(clk), .RSTB(n2266), .Q(\r[11][2] )
         );
  DFFARX1 \r_reg[11][1]  ( .D(n401), .CLK(clk), .RSTB(n2266), .Q(\r[11][1] )
         );
  DFFARX1 \r_reg[11][0]  ( .D(n400), .CLK(clk), .RSTB(n2266), .Q(\r[11][0] )
         );
  DFFARX1 \r_reg[10][31]  ( .D(n399), .CLK(clk), .RSTB(n2267), .Q(\r[10][31] )
         );
  DFFARX1 \r_reg[10][30]  ( .D(n398), .CLK(clk), .RSTB(n2267), .Q(\r[10][30] )
         );
  DFFARX1 \r_reg[10][29]  ( .D(n397), .CLK(clk), .RSTB(n2267), .Q(\r[10][29] )
         );
  DFFARX1 \r_reg[10][28]  ( .D(n396), .CLK(clk), .RSTB(n2267), .Q(\r[10][28] )
         );
  DFFARX1 \r_reg[10][27]  ( .D(n395), .CLK(clk), .RSTB(n2267), .Q(\r[10][27] )
         );
  DFFARX1 \r_reg[10][26]  ( .D(n394), .CLK(clk), .RSTB(n2267), .Q(\r[10][26] )
         );
  DFFARX1 \r_reg[10][25]  ( .D(n393), .CLK(clk), .RSTB(n2267), .Q(\r[10][25] )
         );
  DFFARX1 \r_reg[10][24]  ( .D(n392), .CLK(clk), .RSTB(n2267), .Q(\r[10][24] )
         );
  DFFARX1 \r_reg[10][23]  ( .D(n391), .CLK(clk), .RSTB(n2267), .Q(\r[10][23] )
         );
  DFFARX1 \r_reg[10][22]  ( .D(n390), .CLK(clk), .RSTB(n2267), .Q(\r[10][22] )
         );
  DFFARX1 \r_reg[10][21]  ( .D(n389), .CLK(clk), .RSTB(n2267), .Q(\r[10][21] )
         );
  DFFARX1 \r_reg[10][20]  ( .D(n388), .CLK(clk), .RSTB(n2267), .Q(\r[10][20] )
         );
  DFFARX1 \r_reg[10][19]  ( .D(n387), .CLK(clk), .RSTB(n2268), .Q(\r[10][19] )
         );
  DFFARX1 \r_reg[10][18]  ( .D(n386), .CLK(clk), .RSTB(n2268), .Q(\r[10][18] )
         );
  DFFARX1 \r_reg[10][17]  ( .D(n385), .CLK(clk), .RSTB(n2268), .Q(\r[10][17] )
         );
  DFFARX1 \r_reg[10][16]  ( .D(n384), .CLK(clk), .RSTB(n2268), .Q(\r[10][16] )
         );
  DFFARX1 \r_reg[10][15]  ( .D(n383), .CLK(clk), .RSTB(n2268), .Q(\r[10][15] )
         );
  DFFARX1 \r_reg[10][14]  ( .D(n382), .CLK(clk), .RSTB(n2268), .Q(\r[10][14] )
         );
  DFFARX1 \r_reg[10][13]  ( .D(n381), .CLK(clk), .RSTB(n2268), .Q(\r[10][13] )
         );
  DFFARX1 \r_reg[10][12]  ( .D(n380), .CLK(clk), .RSTB(n2268), .Q(\r[10][12] )
         );
  DFFARX1 \r_reg[10][11]  ( .D(n379), .CLK(clk), .RSTB(n2268), .Q(\r[10][11] )
         );
  DFFARX1 \r_reg[10][10]  ( .D(n378), .CLK(clk), .RSTB(n2268), .Q(\r[10][10] )
         );
  DFFARX1 \r_reg[10][9]  ( .D(n377), .CLK(clk), .RSTB(n2268), .Q(\r[10][9] )
         );
  DFFARX1 \r_reg[10][8]  ( .D(n376), .CLK(clk), .RSTB(n2268), .Q(\r[10][8] )
         );
  DFFARX1 \r_reg[10][7]  ( .D(n375), .CLK(clk), .RSTB(n2269), .Q(\r[10][7] )
         );
  DFFARX1 \r_reg[10][6]  ( .D(n374), .CLK(clk), .RSTB(n2269), .Q(\r[10][6] )
         );
  DFFARX1 \r_reg[10][5]  ( .D(n373), .CLK(clk), .RSTB(n2269), .Q(\r[10][5] )
         );
  DFFARX1 \r_reg[10][4]  ( .D(n372), .CLK(clk), .RSTB(n2269), .Q(\r[10][4] )
         );
  DFFARX1 \r_reg[10][3]  ( .D(n371), .CLK(clk), .RSTB(n2269), .Q(\r[10][3] )
         );
  DFFARX1 \r_reg[10][2]  ( .D(n370), .CLK(clk), .RSTB(n2269), .Q(\r[10][2] )
         );
  DFFARX1 \r_reg[10][1]  ( .D(n369), .CLK(clk), .RSTB(n2269), .Q(\r[10][1] )
         );
  DFFARX1 \r_reg[10][0]  ( .D(n368), .CLK(clk), .RSTB(n2269), .Q(\r[10][0] )
         );
  DFFARX1 \r_reg[9][31]  ( .D(n367), .CLK(clk), .RSTB(n2269), .Q(\r[9][31] )
         );
  DFFARX1 \r_reg[9][30]  ( .D(n366), .CLK(clk), .RSTB(n2269), .Q(\r[9][30] )
         );
  DFFARX1 \r_reg[9][29]  ( .D(n365), .CLK(clk), .RSTB(n2269), .Q(\r[9][29] )
         );
  DFFARX1 \r_reg[9][28]  ( .D(n364), .CLK(clk), .RSTB(n2269), .Q(\r[9][28] )
         );
  DFFARX1 \r_reg[9][27]  ( .D(n363), .CLK(clk), .RSTB(n2270), .Q(\r[9][27] )
         );
  DFFARX1 \r_reg[9][26]  ( .D(n362), .CLK(clk), .RSTB(n2270), .Q(\r[9][26] )
         );
  DFFARX1 \r_reg[9][25]  ( .D(n361), .CLK(clk), .RSTB(n2270), .Q(\r[9][25] )
         );
  DFFARX1 \r_reg[9][24]  ( .D(n360), .CLK(clk), .RSTB(n2270), .Q(\r[9][24] )
         );
  DFFARX1 \r_reg[9][23]  ( .D(n359), .CLK(clk), .RSTB(n2270), .Q(\r[9][23] )
         );
  DFFARX1 \r_reg[9][22]  ( .D(n358), .CLK(clk), .RSTB(n2270), .Q(\r[9][22] )
         );
  DFFARX1 \r_reg[9][21]  ( .D(n357), .CLK(clk), .RSTB(n2270), .Q(\r[9][21] )
         );
  DFFARX1 \r_reg[9][20]  ( .D(n356), .CLK(clk), .RSTB(n2270), .Q(\r[9][20] )
         );
  DFFARX1 \r_reg[9][19]  ( .D(n355), .CLK(clk), .RSTB(n2270), .Q(\r[9][19] )
         );
  DFFARX1 \r_reg[9][18]  ( .D(n354), .CLK(clk), .RSTB(n2270), .Q(\r[9][18] )
         );
  DFFARX1 \r_reg[9][17]  ( .D(n353), .CLK(clk), .RSTB(n2270), .Q(\r[9][17] )
         );
  DFFARX1 \r_reg[9][16]  ( .D(n352), .CLK(clk), .RSTB(n2270), .Q(\r[9][16] )
         );
  DFFARX1 \r_reg[9][15]  ( .D(n351), .CLK(clk), .RSTB(n2271), .Q(\r[9][15] )
         );
  DFFARX1 \r_reg[9][14]  ( .D(n350), .CLK(clk), .RSTB(n2271), .Q(\r[9][14] )
         );
  DFFARX1 \r_reg[9][13]  ( .D(n349), .CLK(clk), .RSTB(n2271), .Q(\r[9][13] )
         );
  DFFARX1 \r_reg[9][12]  ( .D(n348), .CLK(clk), .RSTB(n2271), .Q(\r[9][12] )
         );
  DFFARX1 \r_reg[9][11]  ( .D(n347), .CLK(clk), .RSTB(n2271), .Q(\r[9][11] )
         );
  DFFARX1 \r_reg[9][10]  ( .D(n346), .CLK(clk), .RSTB(n2271), .Q(\r[9][10] )
         );
  DFFARX1 \r_reg[9][9]  ( .D(n345), .CLK(clk), .RSTB(n2271), .Q(\r[9][9] ) );
  DFFARX1 \r_reg[9][8]  ( .D(n344), .CLK(clk), .RSTB(n2271), .Q(\r[9][8] ) );
  DFFARX1 \r_reg[9][7]  ( .D(n343), .CLK(clk), .RSTB(n2271), .Q(\r[9][7] ) );
  DFFARX1 \r_reg[9][6]  ( .D(n342), .CLK(clk), .RSTB(n2271), .Q(\r[9][6] ) );
  DFFARX1 \r_reg[9][5]  ( .D(n341), .CLK(clk), .RSTB(n2271), .Q(\r[9][5] ) );
  DFFARX1 \r_reg[9][4]  ( .D(n340), .CLK(clk), .RSTB(n2271), .Q(\r[9][4] ) );
  DFFARX1 \r_reg[9][3]  ( .D(n339), .CLK(clk), .RSTB(n2272), .Q(\r[9][3] ) );
  DFFARX1 \r_reg[9][2]  ( .D(n338), .CLK(clk), .RSTB(n2272), .Q(\r[9][2] ) );
  DFFARX1 \r_reg[9][1]  ( .D(n337), .CLK(clk), .RSTB(n2272), .Q(\r[9][1] ) );
  DFFARX1 \r_reg[9][0]  ( .D(n336), .CLK(clk), .RSTB(n2272), .Q(\r[9][0] ) );
  DFFARX1 \r_reg[8][31]  ( .D(n335), .CLK(clk), .RSTB(n2272), .Q(\r[8][31] )
         );
  DFFARX1 \r_reg[8][30]  ( .D(n334), .CLK(clk), .RSTB(n2272), .Q(\r[8][30] )
         );
  DFFARX1 \r_reg[8][29]  ( .D(n333), .CLK(clk), .RSTB(n2272), .Q(\r[8][29] )
         );
  DFFARX1 \r_reg[8][28]  ( .D(n332), .CLK(clk), .RSTB(n2272), .Q(\r[8][28] )
         );
  DFFARX1 \r_reg[8][27]  ( .D(n331), .CLK(clk), .RSTB(n2272), .Q(\r[8][27] )
         );
  DFFARX1 \r_reg[8][26]  ( .D(n330), .CLK(clk), .RSTB(n2272), .Q(\r[8][26] )
         );
  DFFARX1 \r_reg[8][25]  ( .D(n329), .CLK(clk), .RSTB(n2272), .Q(\r[8][25] )
         );
  DFFARX1 \r_reg[8][24]  ( .D(n328), .CLK(clk), .RSTB(n2272), .Q(\r[8][24] )
         );
  DFFARX1 \r_reg[8][23]  ( .D(n327), .CLK(clk), .RSTB(n2273), .Q(\r[8][23] )
         );
  DFFARX1 \r_reg[8][22]  ( .D(n326), .CLK(clk), .RSTB(n2273), .Q(\r[8][22] )
         );
  DFFARX1 \r_reg[8][21]  ( .D(n325), .CLK(clk), .RSTB(n2273), .Q(\r[8][21] )
         );
  DFFARX1 \r_reg[8][20]  ( .D(n324), .CLK(clk), .RSTB(n2273), .Q(\r[8][20] )
         );
  DFFARX1 \r_reg[8][19]  ( .D(n323), .CLK(clk), .RSTB(n2273), .Q(\r[8][19] )
         );
  DFFARX1 \r_reg[8][18]  ( .D(n322), .CLK(clk), .RSTB(n2273), .Q(\r[8][18] )
         );
  DFFARX1 \r_reg[8][17]  ( .D(n321), .CLK(clk), .RSTB(n2273), .Q(\r[8][17] )
         );
  DFFARX1 \r_reg[8][16]  ( .D(n320), .CLK(clk), .RSTB(n2273), .Q(\r[8][16] )
         );
  DFFARX1 \r_reg[8][15]  ( .D(n319), .CLK(clk), .RSTB(n2273), .Q(\r[8][15] )
         );
  DFFARX1 \r_reg[8][14]  ( .D(n318), .CLK(clk), .RSTB(n2273), .Q(\r[8][14] )
         );
  DFFARX1 \r_reg[8][13]  ( .D(n317), .CLK(clk), .RSTB(n2273), .Q(\r[8][13] )
         );
  DFFARX1 \r_reg[8][12]  ( .D(n316), .CLK(clk), .RSTB(n2273), .Q(\r[8][12] )
         );
  DFFARX1 \r_reg[8][11]  ( .D(n315), .CLK(clk), .RSTB(n2274), .Q(\r[8][11] )
         );
  DFFARX1 \r_reg[8][10]  ( .D(n314), .CLK(clk), .RSTB(n2274), .Q(\r[8][10] )
         );
  DFFARX1 \r_reg[8][9]  ( .D(n313), .CLK(clk), .RSTB(n2274), .Q(\r[8][9] ) );
  DFFARX1 \r_reg[8][8]  ( .D(n312), .CLK(clk), .RSTB(n2274), .Q(\r[8][8] ) );
  DFFARX1 \r_reg[8][7]  ( .D(n311), .CLK(clk), .RSTB(n2274), .Q(\r[8][7] ) );
  DFFARX1 \r_reg[8][6]  ( .D(n310), .CLK(clk), .RSTB(n2274), .Q(\r[8][6] ) );
  DFFARX1 \r_reg[8][5]  ( .D(n309), .CLK(clk), .RSTB(n2274), .Q(\r[8][5] ) );
  DFFARX1 \r_reg[8][4]  ( .D(n308), .CLK(clk), .RSTB(n2274), .Q(\r[8][4] ) );
  DFFARX1 \r_reg[8][3]  ( .D(n307), .CLK(clk), .RSTB(n2274), .Q(\r[8][3] ) );
  DFFARX1 \r_reg[8][2]  ( .D(n306), .CLK(clk), .RSTB(n2274), .Q(\r[8][2] ) );
  DFFARX1 \r_reg[8][1]  ( .D(n305), .CLK(clk), .RSTB(n2274), .Q(\r[8][1] ) );
  DFFARX1 \r_reg[8][0]  ( .D(n304), .CLK(clk), .RSTB(n2274), .Q(\r[8][0] ) );
  DFFARX1 \r_reg[7][31]  ( .D(n303), .CLK(clk), .RSTB(n2275), .Q(\r[7][31] )
         );
  DFFARX1 \r_reg[7][30]  ( .D(n302), .CLK(clk), .RSTB(n2275), .Q(\r[7][30] )
         );
  DFFARX1 \r_reg[7][29]  ( .D(n301), .CLK(clk), .RSTB(n2275), .Q(\r[7][29] )
         );
  DFFARX1 \r_reg[7][28]  ( .D(n300), .CLK(clk), .RSTB(n2275), .Q(\r[7][28] )
         );
  DFFARX1 \r_reg[7][27]  ( .D(n299), .CLK(clk), .RSTB(n2275), .Q(\r[7][27] )
         );
  DFFARX1 \r_reg[7][26]  ( .D(n298), .CLK(clk), .RSTB(n2275), .Q(\r[7][26] )
         );
  DFFARX1 \r_reg[7][25]  ( .D(n297), .CLK(clk), .RSTB(n2275), .Q(\r[7][25] )
         );
  DFFARX1 \r_reg[7][24]  ( .D(n296), .CLK(clk), .RSTB(n2275), .Q(\r[7][24] )
         );
  DFFARX1 \r_reg[7][23]  ( .D(n295), .CLK(clk), .RSTB(n2275), .Q(\r[7][23] )
         );
  DFFARX1 \r_reg[7][22]  ( .D(n294), .CLK(clk), .RSTB(n2275), .Q(\r[7][22] )
         );
  DFFARX1 \r_reg[7][21]  ( .D(n293), .CLK(clk), .RSTB(n2275), .Q(\r[7][21] )
         );
  DFFARX1 \r_reg[7][20]  ( .D(n292), .CLK(clk), .RSTB(n2275), .Q(\r[7][20] )
         );
  DFFARX1 \r_reg[7][19]  ( .D(n291), .CLK(clk), .RSTB(n2276), .Q(\r[7][19] )
         );
  DFFARX1 \r_reg[7][18]  ( .D(n290), .CLK(clk), .RSTB(n2276), .Q(\r[7][18] )
         );
  DFFARX1 \r_reg[7][17]  ( .D(n289), .CLK(clk), .RSTB(n2276), .Q(\r[7][17] )
         );
  DFFARX1 \r_reg[7][16]  ( .D(n288), .CLK(clk), .RSTB(n2276), .Q(\r[7][16] )
         );
  DFFARX1 \r_reg[7][15]  ( .D(n287), .CLK(clk), .RSTB(n2276), .Q(\r[7][15] )
         );
  DFFARX1 \r_reg[7][14]  ( .D(n286), .CLK(clk), .RSTB(n2276), .Q(\r[7][14] )
         );
  DFFARX1 \r_reg[7][13]  ( .D(n285), .CLK(clk), .RSTB(n2276), .Q(\r[7][13] )
         );
  DFFARX1 \r_reg[7][12]  ( .D(n284), .CLK(clk), .RSTB(n2276), .Q(\r[7][12] )
         );
  DFFARX1 \r_reg[7][11]  ( .D(n283), .CLK(clk), .RSTB(n2276), .Q(\r[7][11] )
         );
  DFFARX1 \r_reg[7][10]  ( .D(n282), .CLK(clk), .RSTB(n2276), .Q(\r[7][10] )
         );
  DFFARX1 \r_reg[7][9]  ( .D(n281), .CLK(clk), .RSTB(n2276), .Q(\r[7][9] ) );
  DFFARX1 \r_reg[7][8]  ( .D(n280), .CLK(clk), .RSTB(n2276), .Q(\r[7][8] ) );
  DFFARX1 \r_reg[7][7]  ( .D(n279), .CLK(clk), .RSTB(n2277), .Q(\r[7][7] ) );
  DFFARX1 \r_reg[7][6]  ( .D(n278), .CLK(clk), .RSTB(n2277), .Q(\r[7][6] ) );
  DFFARX1 \r_reg[7][5]  ( .D(n277), .CLK(clk), .RSTB(n2277), .Q(\r[7][5] ) );
  DFFARX1 \r_reg[7][4]  ( .D(n276), .CLK(clk), .RSTB(n2277), .Q(\r[7][4] ) );
  DFFARX1 \r_reg[7][3]  ( .D(n275), .CLK(clk), .RSTB(n2277), .Q(\r[7][3] ) );
  DFFARX1 \r_reg[7][2]  ( .D(n274), .CLK(clk), .RSTB(n2277), .Q(\r[7][2] ) );
  DFFARX1 \r_reg[7][1]  ( .D(n273), .CLK(clk), .RSTB(n2277), .Q(\r[7][1] ) );
  DFFARX1 \r_reg[7][0]  ( .D(n272), .CLK(clk), .RSTB(n2277), .Q(\r[7][0] ) );
  DFFARX1 \r_reg[6][31]  ( .D(n271), .CLK(clk), .RSTB(n2277), .Q(\r[6][31] )
         );
  DFFARX1 \r_reg[6][30]  ( .D(n270), .CLK(clk), .RSTB(n2277), .Q(\r[6][30] )
         );
  DFFARX1 \r_reg[6][29]  ( .D(n269), .CLK(clk), .RSTB(n2277), .Q(\r[6][29] )
         );
  DFFARX1 \r_reg[6][28]  ( .D(n268), .CLK(clk), .RSTB(n2277), .Q(\r[6][28] )
         );
  DFFARX1 \r_reg[6][27]  ( .D(n267), .CLK(clk), .RSTB(n2278), .Q(\r[6][27] )
         );
  DFFARX1 \r_reg[6][26]  ( .D(n266), .CLK(clk), .RSTB(n2278), .Q(\r[6][26] )
         );
  DFFARX1 \r_reg[6][25]  ( .D(n265), .CLK(clk), .RSTB(n2278), .Q(\r[6][25] )
         );
  DFFARX1 \r_reg[6][24]  ( .D(n264), .CLK(clk), .RSTB(n2278), .Q(\r[6][24] )
         );
  DFFARX1 \r_reg[6][23]  ( .D(n263), .CLK(clk), .RSTB(n2278), .Q(\r[6][23] )
         );
  DFFARX1 \r_reg[6][22]  ( .D(n262), .CLK(clk), .RSTB(n2278), .Q(\r[6][22] )
         );
  DFFARX1 \r_reg[6][21]  ( .D(n261), .CLK(clk), .RSTB(n2278), .Q(\r[6][21] )
         );
  DFFARX1 \r_reg[6][20]  ( .D(n260), .CLK(clk), .RSTB(n2278), .Q(\r[6][20] )
         );
  DFFARX1 \r_reg[6][19]  ( .D(n259), .CLK(clk), .RSTB(n2278), .Q(\r[6][19] )
         );
  DFFARX1 \r_reg[6][18]  ( .D(n258), .CLK(clk), .RSTB(n2278), .Q(\r[6][18] )
         );
  DFFARX1 \r_reg[6][17]  ( .D(n257), .CLK(clk), .RSTB(n2278), .Q(\r[6][17] )
         );
  DFFARX1 \r_reg[6][16]  ( .D(n256), .CLK(clk), .RSTB(n2278), .Q(\r[6][16] )
         );
  DFFARX1 \r_reg[6][15]  ( .D(n255), .CLK(clk), .RSTB(n2279), .Q(\r[6][15] )
         );
  DFFARX1 \r_reg[6][14]  ( .D(n254), .CLK(clk), .RSTB(n2279), .Q(\r[6][14] )
         );
  DFFARX1 \r_reg[6][13]  ( .D(n253), .CLK(clk), .RSTB(n2279), .Q(\r[6][13] )
         );
  DFFARX1 \r_reg[6][12]  ( .D(n252), .CLK(clk), .RSTB(n2279), .Q(\r[6][12] )
         );
  DFFARX1 \r_reg[6][11]  ( .D(n251), .CLK(clk), .RSTB(n2279), .Q(\r[6][11] )
         );
  DFFARX1 \r_reg[6][10]  ( .D(n250), .CLK(clk), .RSTB(n2279), .Q(\r[6][10] )
         );
  DFFARX1 \r_reg[6][9]  ( .D(n249), .CLK(clk), .RSTB(n2279), .Q(\r[6][9] ) );
  DFFARX1 \r_reg[6][8]  ( .D(n248), .CLK(clk), .RSTB(n2279), .Q(\r[6][8] ) );
  DFFARX1 \r_reg[6][7]  ( .D(n247), .CLK(clk), .RSTB(n2279), .Q(\r[6][7] ) );
  DFFARX1 \r_reg[6][6]  ( .D(n246), .CLK(clk), .RSTB(n2279), .Q(\r[6][6] ) );
  DFFARX1 \r_reg[6][5]  ( .D(n245), .CLK(clk), .RSTB(n2279), .Q(\r[6][5] ) );
  DFFARX1 \r_reg[6][4]  ( .D(n244), .CLK(clk), .RSTB(n2279), .Q(\r[6][4] ) );
  DFFARX1 \r_reg[6][3]  ( .D(n243), .CLK(clk), .RSTB(n2280), .Q(\r[6][3] ) );
  DFFARX1 \r_reg[6][2]  ( .D(n242), .CLK(clk), .RSTB(n2280), .Q(\r[6][2] ) );
  DFFARX1 \r_reg[6][1]  ( .D(n241), .CLK(clk), .RSTB(n2280), .Q(\r[6][1] ) );
  DFFARX1 \r_reg[6][0]  ( .D(n240), .CLK(clk), .RSTB(n2280), .Q(\r[6][0] ) );
  DFFARX1 \r_reg[5][31]  ( .D(n239), .CLK(clk), .RSTB(n2280), .Q(\r[5][31] )
         );
  DFFARX1 \r_reg[5][30]  ( .D(n238), .CLK(clk), .RSTB(n2280), .Q(\r[5][30] )
         );
  DFFARX1 \r_reg[5][29]  ( .D(n237), .CLK(clk), .RSTB(n2280), .Q(\r[5][29] )
         );
  DFFARX1 \r_reg[5][28]  ( .D(n236), .CLK(clk), .RSTB(n2280), .Q(\r[5][28] )
         );
  DFFARX1 \r_reg[5][27]  ( .D(n235), .CLK(clk), .RSTB(n2280), .Q(\r[5][27] )
         );
  DFFARX1 \r_reg[5][26]  ( .D(n234), .CLK(clk), .RSTB(n2280), .Q(\r[5][26] )
         );
  DFFARX1 \r_reg[5][25]  ( .D(n233), .CLK(clk), .RSTB(n2280), .Q(\r[5][25] )
         );
  DFFARX1 \r_reg[5][24]  ( .D(n232), .CLK(clk), .RSTB(n2280), .Q(\r[5][24] )
         );
  DFFARX1 \r_reg[5][23]  ( .D(n231), .CLK(clk), .RSTB(n2281), .Q(\r[5][23] )
         );
  DFFARX1 \r_reg[5][22]  ( .D(n230), .CLK(clk), .RSTB(n2281), .Q(\r[5][22] )
         );
  DFFARX1 \r_reg[5][21]  ( .D(n229), .CLK(clk), .RSTB(n2281), .Q(\r[5][21] )
         );
  DFFARX1 \r_reg[5][20]  ( .D(n228), .CLK(clk), .RSTB(n2281), .Q(\r[5][20] )
         );
  DFFARX1 \r_reg[5][19]  ( .D(n227), .CLK(clk), .RSTB(n2281), .Q(\r[5][19] )
         );
  DFFARX1 \r_reg[5][18]  ( .D(n226), .CLK(clk), .RSTB(n2281), .Q(\r[5][18] )
         );
  DFFARX1 \r_reg[5][17]  ( .D(n225), .CLK(clk), .RSTB(n2281), .Q(\r[5][17] )
         );
  DFFARX1 \r_reg[5][16]  ( .D(n224), .CLK(clk), .RSTB(n2281), .Q(\r[5][16] )
         );
  DFFARX1 \r_reg[5][15]  ( .D(n223), .CLK(clk), .RSTB(n2281), .Q(\r[5][15] )
         );
  DFFARX1 \r_reg[5][14]  ( .D(n222), .CLK(clk), .RSTB(n2281), .Q(\r[5][14] )
         );
  DFFARX1 \r_reg[5][13]  ( .D(n221), .CLK(clk), .RSTB(n2281), .Q(\r[5][13] )
         );
  DFFARX1 \r_reg[5][12]  ( .D(n220), .CLK(clk), .RSTB(n2281), .Q(\r[5][12] )
         );
  DFFARX1 \r_reg[5][11]  ( .D(n219), .CLK(clk), .RSTB(n2282), .Q(\r[5][11] )
         );
  DFFARX1 \r_reg[5][10]  ( .D(n218), .CLK(clk), .RSTB(n2282), .Q(\r[5][10] )
         );
  DFFARX1 \r_reg[5][9]  ( .D(n217), .CLK(clk), .RSTB(n2282), .Q(\r[5][9] ) );
  DFFARX1 \r_reg[5][8]  ( .D(n216), .CLK(clk), .RSTB(n2282), .Q(\r[5][8] ) );
  DFFARX1 \r_reg[5][7]  ( .D(n215), .CLK(clk), .RSTB(n2282), .Q(\r[5][7] ) );
  DFFARX1 \r_reg[5][6]  ( .D(n214), .CLK(clk), .RSTB(n2282), .Q(\r[5][6] ) );
  DFFARX1 \r_reg[5][5]  ( .D(n213), .CLK(clk), .RSTB(n2282), .Q(\r[5][5] ) );
  DFFARX1 \r_reg[5][4]  ( .D(n212), .CLK(clk), .RSTB(n2282), .Q(\r[5][4] ) );
  DFFARX1 \r_reg[5][3]  ( .D(n211), .CLK(clk), .RSTB(n2282), .Q(\r[5][3] ) );
  DFFARX1 \r_reg[5][2]  ( .D(n210), .CLK(clk), .RSTB(n2282), .Q(\r[5][2] ) );
  DFFARX1 \r_reg[5][1]  ( .D(n209), .CLK(clk), .RSTB(n2282), .Q(\r[5][1] ) );
  DFFARX1 \r_reg[5][0]  ( .D(n208), .CLK(clk), .RSTB(n2282), .Q(\r[5][0] ) );
  DFFARX1 \r_reg[4][31]  ( .D(n207), .CLK(clk), .RSTB(n2283), .Q(\r[4][31] )
         );
  DFFARX1 \r_reg[4][30]  ( .D(n206), .CLK(clk), .RSTB(n2283), .Q(\r[4][30] )
         );
  DFFARX1 \r_reg[4][29]  ( .D(n205), .CLK(clk), .RSTB(n2283), .Q(\r[4][29] )
         );
  DFFARX1 \r_reg[4][28]  ( .D(n204), .CLK(clk), .RSTB(n2283), .Q(\r[4][28] )
         );
  DFFARX1 \r_reg[4][27]  ( .D(n203), .CLK(clk), .RSTB(n2283), .Q(\r[4][27] )
         );
  DFFARX1 \r_reg[4][26]  ( .D(n202), .CLK(clk), .RSTB(n2283), .Q(\r[4][26] )
         );
  DFFARX1 \r_reg[4][25]  ( .D(n201), .CLK(clk), .RSTB(n2283), .Q(\r[4][25] )
         );
  DFFARX1 \r_reg[4][24]  ( .D(n200), .CLK(clk), .RSTB(n2283), .Q(\r[4][24] )
         );
  DFFARX1 \r_reg[4][23]  ( .D(n199), .CLK(clk), .RSTB(n2283), .Q(\r[4][23] )
         );
  DFFARX1 \r_reg[4][22]  ( .D(n198), .CLK(clk), .RSTB(n2283), .Q(\r[4][22] )
         );
  DFFARX1 \r_reg[4][21]  ( .D(n197), .CLK(clk), .RSTB(n2283), .Q(\r[4][21] )
         );
  DFFARX1 \r_reg[4][20]  ( .D(n196), .CLK(clk), .RSTB(n2283), .Q(\r[4][20] )
         );
  DFFARX1 \r_reg[4][19]  ( .D(n195), .CLK(clk), .RSTB(n2284), .Q(\r[4][19] )
         );
  DFFARX1 \r_reg[4][18]  ( .D(n194), .CLK(clk), .RSTB(n2284), .Q(\r[4][18] )
         );
  DFFARX1 \r_reg[4][17]  ( .D(n193), .CLK(clk), .RSTB(n2284), .Q(\r[4][17] )
         );
  DFFARX1 \r_reg[4][16]  ( .D(n192), .CLK(clk), .RSTB(n2284), .Q(\r[4][16] )
         );
  DFFARX1 \r_reg[4][15]  ( .D(n191), .CLK(clk), .RSTB(n2284), .Q(\r[4][15] )
         );
  DFFARX1 \r_reg[4][14]  ( .D(n190), .CLK(clk), .RSTB(n2284), .Q(\r[4][14] )
         );
  DFFARX1 \r_reg[4][13]  ( .D(n189), .CLK(clk), .RSTB(n2284), .Q(\r[4][13] )
         );
  DFFARX1 \r_reg[4][12]  ( .D(n188), .CLK(clk), .RSTB(n2284), .Q(\r[4][12] )
         );
  DFFARX1 \r_reg[4][11]  ( .D(n187), .CLK(clk), .RSTB(n2284), .Q(\r[4][11] )
         );
  DFFARX1 \r_reg[4][10]  ( .D(n186), .CLK(clk), .RSTB(n2284), .Q(\r[4][10] )
         );
  DFFARX1 \r_reg[4][9]  ( .D(n185), .CLK(clk), .RSTB(n2284), .Q(\r[4][9] ) );
  DFFARX1 \r_reg[4][8]  ( .D(n184), .CLK(clk), .RSTB(n2284), .Q(\r[4][8] ) );
  DFFARX1 \r_reg[4][7]  ( .D(n183), .CLK(clk), .RSTB(n2285), .Q(\r[4][7] ) );
  DFFARX1 \r_reg[4][6]  ( .D(n182), .CLK(clk), .RSTB(n2285), .Q(\r[4][6] ) );
  DFFARX1 \r_reg[4][5]  ( .D(n181), .CLK(clk), .RSTB(n2285), .Q(\r[4][5] ) );
  DFFARX1 \r_reg[4][4]  ( .D(n180), .CLK(clk), .RSTB(n2285), .Q(\r[4][4] ) );
  DFFARX1 \r_reg[4][3]  ( .D(n179), .CLK(clk), .RSTB(n2285), .Q(\r[4][3] ) );
  DFFARX1 \r_reg[4][2]  ( .D(n178), .CLK(clk), .RSTB(n2285), .Q(\r[4][2] ) );
  DFFARX1 \r_reg[4][1]  ( .D(n177), .CLK(clk), .RSTB(n2285), .Q(\r[4][1] ) );
  DFFARX1 \r_reg[4][0]  ( .D(n176), .CLK(clk), .RSTB(n2285), .Q(\r[4][0] ) );
  DFFARX1 \r_reg[3][31]  ( .D(n175), .CLK(clk), .RSTB(n2285), .Q(\r[3][31] )
         );
  DFFARX1 \r_reg[3][30]  ( .D(n174), .CLK(clk), .RSTB(n2285), .Q(\r[3][30] )
         );
  DFFARX1 \r_reg[3][29]  ( .D(n173), .CLK(clk), .RSTB(n2285), .Q(\r[3][29] )
         );
  DFFARX1 \r_reg[3][28]  ( .D(n172), .CLK(clk), .RSTB(n2285), .Q(\r[3][28] )
         );
  DFFARX1 \r_reg[3][27]  ( .D(n171), .CLK(clk), .RSTB(n2286), .Q(\r[3][27] )
         );
  DFFARX1 \r_reg[3][26]  ( .D(n170), .CLK(clk), .RSTB(n2286), .Q(\r[3][26] )
         );
  DFFARX1 \r_reg[3][25]  ( .D(n169), .CLK(clk), .RSTB(n2286), .Q(\r[3][25] )
         );
  DFFARX1 \r_reg[3][24]  ( .D(n168), .CLK(clk), .RSTB(n2286), .Q(\r[3][24] )
         );
  DFFARX1 \r_reg[3][23]  ( .D(n167), .CLK(clk), .RSTB(n2286), .Q(\r[3][23] )
         );
  DFFARX1 \r_reg[3][22]  ( .D(n166), .CLK(clk), .RSTB(n2286), .Q(\r[3][22] )
         );
  DFFARX1 \r_reg[3][21]  ( .D(n165), .CLK(clk), .RSTB(n2286), .Q(\r[3][21] )
         );
  DFFARX1 \r_reg[3][20]  ( .D(n164), .CLK(clk), .RSTB(n2286), .Q(\r[3][20] )
         );
  DFFARX1 \r_reg[3][19]  ( .D(n163), .CLK(clk), .RSTB(n2286), .Q(\r[3][19] )
         );
  DFFARX1 \r_reg[3][18]  ( .D(n162), .CLK(clk), .RSTB(n2286), .Q(\r[3][18] )
         );
  DFFARX1 \r_reg[3][17]  ( .D(n161), .CLK(clk), .RSTB(n2286), .Q(\r[3][17] )
         );
  DFFARX1 \r_reg[3][16]  ( .D(n160), .CLK(clk), .RSTB(n2286), .Q(\r[3][16] )
         );
  DFFARX1 \r_reg[3][15]  ( .D(n159), .CLK(clk), .RSTB(n2287), .Q(\r[3][15] )
         );
  DFFARX1 \r_reg[3][14]  ( .D(n158), .CLK(clk), .RSTB(n2287), .Q(\r[3][14] )
         );
  DFFARX1 \r_reg[3][13]  ( .D(n157), .CLK(clk), .RSTB(n2287), .Q(\r[3][13] )
         );
  DFFARX1 \r_reg[3][12]  ( .D(n156), .CLK(clk), .RSTB(n2287), .Q(\r[3][12] )
         );
  DFFARX1 \r_reg[3][11]  ( .D(n155), .CLK(clk), .RSTB(n2287), .Q(\r[3][11] )
         );
  DFFARX1 \r_reg[3][10]  ( .D(n154), .CLK(clk), .RSTB(n2287), .Q(\r[3][10] )
         );
  DFFARX1 \r_reg[3][9]  ( .D(n153), .CLK(clk), .RSTB(n2287), .Q(\r[3][9] ) );
  DFFARX1 \r_reg[3][8]  ( .D(n152), .CLK(clk), .RSTB(n2287), .Q(\r[3][8] ) );
  DFFARX1 \r_reg[3][7]  ( .D(n151), .CLK(clk), .RSTB(n2287), .Q(\r[3][7] ) );
  DFFARX1 \r_reg[3][6]  ( .D(n150), .CLK(clk), .RSTB(n2287), .Q(\r[3][6] ) );
  DFFARX1 \r_reg[3][5]  ( .D(n149), .CLK(clk), .RSTB(n2287), .Q(\r[3][5] ) );
  DFFARX1 \r_reg[3][4]  ( .D(n148), .CLK(clk), .RSTB(n2287), .Q(\r[3][4] ) );
  DFFARX1 \r_reg[3][3]  ( .D(n147), .CLK(clk), .RSTB(n2288), .Q(\r[3][3] ) );
  DFFARX1 \r_reg[3][2]  ( .D(n146), .CLK(clk), .RSTB(n2288), .Q(\r[3][2] ) );
  DFFARX1 \r_reg[3][1]  ( .D(n145), .CLK(clk), .RSTB(n2288), .Q(\r[3][1] ) );
  DFFARX1 \r_reg[3][0]  ( .D(n144), .CLK(clk), .RSTB(n2288), .Q(\r[3][0] ) );
  DFFARX1 \r_reg[2][31]  ( .D(n143), .CLK(clk), .RSTB(n2288), .Q(\r[2][31] )
         );
  DFFARX1 \r_reg[2][30]  ( .D(n142), .CLK(clk), .RSTB(n2288), .Q(\r[2][30] )
         );
  DFFARX1 \r_reg[2][29]  ( .D(n141), .CLK(clk), .RSTB(n2288), .Q(\r[2][29] )
         );
  DFFARX1 \r_reg[2][28]  ( .D(n140), .CLK(clk), .RSTB(n2288), .Q(\r[2][28] )
         );
  DFFARX1 \r_reg[2][27]  ( .D(n139), .CLK(clk), .RSTB(n2288), .Q(\r[2][27] )
         );
  DFFARX1 \r_reg[2][26]  ( .D(n138), .CLK(clk), .RSTB(n2288), .Q(\r[2][26] )
         );
  DFFARX1 \r_reg[2][25]  ( .D(n137), .CLK(clk), .RSTB(n2288), .Q(\r[2][25] )
         );
  DFFARX1 \r_reg[2][24]  ( .D(n136), .CLK(clk), .RSTB(n2288), .Q(\r[2][24] )
         );
  DFFARX1 \r_reg[2][23]  ( .D(n135), .CLK(clk), .RSTB(n2289), .Q(\r[2][23] )
         );
  DFFARX1 \r_reg[2][22]  ( .D(n134), .CLK(clk), .RSTB(n2289), .Q(\r[2][22] )
         );
  DFFARX1 \r_reg[2][21]  ( .D(n133), .CLK(clk), .RSTB(n2289), .Q(\r[2][21] )
         );
  DFFARX1 \r_reg[2][20]  ( .D(n132), .CLK(clk), .RSTB(n2289), .Q(\r[2][20] )
         );
  DFFARX1 \r_reg[2][19]  ( .D(n131), .CLK(clk), .RSTB(n2289), .Q(\r[2][19] )
         );
  DFFARX1 \r_reg[2][18]  ( .D(n130), .CLK(clk), .RSTB(n2289), .Q(\r[2][18] )
         );
  DFFARX1 \r_reg[2][17]  ( .D(n129), .CLK(clk), .RSTB(n2289), .Q(\r[2][17] )
         );
  DFFARX1 \r_reg[2][16]  ( .D(n128), .CLK(clk), .RSTB(n2289), .Q(\r[2][16] )
         );
  DFFARX1 \r_reg[2][15]  ( .D(n127), .CLK(clk), .RSTB(n2289), .Q(\r[2][15] )
         );
  DFFARX1 \r_reg[2][14]  ( .D(n126), .CLK(clk), .RSTB(n2289), .Q(\r[2][14] )
         );
  DFFARX1 \r_reg[2][13]  ( .D(n125), .CLK(clk), .RSTB(n2289), .Q(\r[2][13] )
         );
  DFFARX1 \r_reg[2][12]  ( .D(n124), .CLK(clk), .RSTB(n2289), .Q(\r[2][12] )
         );
  DFFARX1 \r_reg[2][11]  ( .D(n123), .CLK(clk), .RSTB(n2290), .Q(\r[2][11] )
         );
  DFFARX1 \r_reg[2][10]  ( .D(n122), .CLK(clk), .RSTB(n2290), .Q(\r[2][10] )
         );
  DFFARX1 \r_reg[2][9]  ( .D(n121), .CLK(clk), .RSTB(n2290), .Q(\r[2][9] ) );
  DFFARX1 \r_reg[2][8]  ( .D(n120), .CLK(clk), .RSTB(n2290), .Q(\r[2][8] ) );
  DFFARX1 \r_reg[2][7]  ( .D(n119), .CLK(clk), .RSTB(n2290), .Q(\r[2][7] ) );
  DFFARX1 \r_reg[2][6]  ( .D(n118), .CLK(clk), .RSTB(n2290), .Q(\r[2][6] ) );
  DFFARX1 \r_reg[2][5]  ( .D(n117), .CLK(clk), .RSTB(n2290), .Q(\r[2][5] ) );
  DFFARX1 \r_reg[2][4]  ( .D(n116), .CLK(clk), .RSTB(n2290), .Q(\r[2][4] ) );
  DFFARX1 \r_reg[2][3]  ( .D(n115), .CLK(clk), .RSTB(n2290), .Q(\r[2][3] ) );
  DFFARX1 \r_reg[2][2]  ( .D(n114), .CLK(clk), .RSTB(n2290), .Q(\r[2][2] ) );
  DFFARX1 \r_reg[2][1]  ( .D(n113), .CLK(clk), .RSTB(n2290), .Q(\r[2][1] ) );
  DFFARX1 \r_reg[2][0]  ( .D(n112), .CLK(clk), .RSTB(n2290), .Q(\r[2][0] ) );
  DFFARX1 \r_reg[1][31]  ( .D(n111), .CLK(clk), .RSTB(n2291), .Q(\r[1][31] )
         );
  DFFARX1 \r_reg[1][30]  ( .D(n110), .CLK(clk), .RSTB(n2291), .Q(\r[1][30] )
         );
  DFFARX1 \r_reg[1][29]  ( .D(n109), .CLK(clk), .RSTB(n2291), .Q(\r[1][29] )
         );
  DFFARX1 \r_reg[1][28]  ( .D(n108), .CLK(clk), .RSTB(n2291), .Q(\r[1][28] )
         );
  DFFARX1 \r_reg[1][27]  ( .D(n107), .CLK(clk), .RSTB(n2291), .Q(\r[1][27] )
         );
  DFFARX1 \r_reg[1][26]  ( .D(n106), .CLK(clk), .RSTB(n2291), .Q(\r[1][26] )
         );
  DFFARX1 \r_reg[1][25]  ( .D(n105), .CLK(clk), .RSTB(n2291), .Q(\r[1][25] )
         );
  DFFARX1 \r_reg[1][24]  ( .D(n104), .CLK(clk), .RSTB(n2291), .Q(\r[1][24] )
         );
  DFFARX1 \r_reg[1][23]  ( .D(n103), .CLK(clk), .RSTB(n2291), .Q(\r[1][23] )
         );
  DFFARX1 \r_reg[1][22]  ( .D(n102), .CLK(clk), .RSTB(n2291), .Q(\r[1][22] )
         );
  DFFARX1 \r_reg[1][21]  ( .D(n101), .CLK(clk), .RSTB(n2291), .Q(\r[1][21] )
         );
  DFFARX1 \r_reg[1][20]  ( .D(n100), .CLK(clk), .RSTB(n2291), .Q(\r[1][20] )
         );
  DFFARX1 \r_reg[1][19]  ( .D(n99), .CLK(clk), .RSTB(n2292), .Q(\r[1][19] ) );
  DFFARX1 \r_reg[1][18]  ( .D(n98), .CLK(clk), .RSTB(n2292), .Q(\r[1][18] ) );
  DFFARX1 \r_reg[1][17]  ( .D(n97), .CLK(clk), .RSTB(n2292), .Q(\r[1][17] ) );
  DFFARX1 \r_reg[1][16]  ( .D(n96), .CLK(clk), .RSTB(n2292), .Q(\r[1][16] ) );
  DFFARX1 \r_reg[1][15]  ( .D(n95), .CLK(clk), .RSTB(n2292), .Q(\r[1][15] ) );
  DFFARX1 \r_reg[1][14]  ( .D(n94), .CLK(clk), .RSTB(n2292), .Q(\r[1][14] ) );
  DFFARX1 \r_reg[1][13]  ( .D(n93), .CLK(clk), .RSTB(n2292), .Q(\r[1][13] ) );
  DFFARX1 \r_reg[1][12]  ( .D(n92), .CLK(clk), .RSTB(n2292), .Q(\r[1][12] ) );
  DFFARX1 \r_reg[1][11]  ( .D(n91), .CLK(clk), .RSTB(n2292), .Q(\r[1][11] ) );
  DFFARX1 \r_reg[1][10]  ( .D(n90), .CLK(clk), .RSTB(n2292), .Q(\r[1][10] ) );
  DFFARX1 \r_reg[1][9]  ( .D(n89), .CLK(clk), .RSTB(n2292), .Q(\r[1][9] ) );
  DFFARX1 \r_reg[1][8]  ( .D(n88), .CLK(clk), .RSTB(n2292), .Q(\r[1][8] ) );
  DFFARX1 \r_reg[1][7]  ( .D(n87), .CLK(clk), .RSTB(nrst), .Q(\r[1][7] ) );
  DFFARX1 \r_reg[1][6]  ( .D(n86), .CLK(clk), .RSTB(nrst), .Q(\r[1][6] ) );
  DFFARX1 \r_reg[1][5]  ( .D(n85), .CLK(clk), .RSTB(nrst), .Q(\r[1][5] ) );
  DFFARX1 \r_reg[1][4]  ( .D(n84), .CLK(clk), .RSTB(nrst), .Q(\r[1][4] ) );
  DFFARX1 \r_reg[1][3]  ( .D(n83), .CLK(clk), .RSTB(nrst), .Q(\r[1][3] ) );
  DFFARX1 \r_reg[1][2]  ( .D(n82), .CLK(clk), .RSTB(nrst), .Q(\r[1][2] ) );
  DFFARX1 \r_reg[1][1]  ( .D(n81), .CLK(clk), .RSTB(nrst), .Q(\r[1][1] ) );
  DFFARX1 \r_reg[1][0]  ( .D(n80), .CLK(clk), .RSTB(nrst), .Q(\r[1][0] ) );
  AO22X1 U101 ( .IN1(wr_data[0]), .IN2(n2208), .IN3(\r[1][0] ), .IN4(n37), .Q(
        n80) );
  AO22X1 U102 ( .IN1(wr_data[1]), .IN2(n2208), .IN3(\r[1][1] ), .IN4(n37), .Q(
        n81) );
  AO22X1 U103 ( .IN1(wr_data[2]), .IN2(n2208), .IN3(\r[1][2] ), .IN4(n37), .Q(
        n82) );
  AO22X1 U104 ( .IN1(wr_data[3]), .IN2(n2208), .IN3(\r[1][3] ), .IN4(n37), .Q(
        n83) );
  AO22X1 U105 ( .IN1(wr_data[4]), .IN2(n2208), .IN3(\r[1][4] ), .IN4(n37), .Q(
        n84) );
  AO22X1 U106 ( .IN1(wr_data[5]), .IN2(n2208), .IN3(\r[1][5] ), .IN4(n37), .Q(
        n85) );
  AO22X1 U107 ( .IN1(wr_data[6]), .IN2(n2208), .IN3(\r[1][6] ), .IN4(n37), .Q(
        n86) );
  AO22X1 U108 ( .IN1(wr_data[7]), .IN2(n2208), .IN3(\r[1][7] ), .IN4(n37), .Q(
        n87) );
  AO22X1 U109 ( .IN1(wr_data[8]), .IN2(n2208), .IN3(\r[1][8] ), .IN4(n2207),
        .Q(n88) );
  AO22X1 U110 ( .IN1(wr_data[9]), .IN2(n2208), .IN3(\r[1][9] ), .IN4(n2207),
        .Q(n89) );
  AO22X1 U111 ( .IN1(wr_data[10]), .IN2(n2209), .IN3(\r[1][10] ), .IN4(n2207),
        .Q(n90) );
  AO22X1 U112 ( .IN1(wr_data[11]), .IN2(n2209), .IN3(\r[1][11] ), .IN4(n2207),
        .Q(n91) );
  AO22X1 U113 ( .IN1(wr_data[12]), .IN2(n2209), .IN3(\r[1][12] ), .IN4(n2207),
        .Q(n92) );
  AO22X1 U114 ( .IN1(wr_data[13]), .IN2(n2209), .IN3(\r[1][13] ), .IN4(n2207),
        .Q(n93) );
  AO22X1 U115 ( .IN1(wr_data[14]), .IN2(n2209), .IN3(\r[1][14] ), .IN4(n2207),
        .Q(n94) );
  AO22X1 U116 ( .IN1(wr_data[15]), .IN2(n2209), .IN3(\r[1][15] ), .IN4(n2207),
        .Q(n95) );
  AO22X1 U117 ( .IN1(wr_data[16]), .IN2(n2209), .IN3(\r[1][16] ), .IN4(n2207),
        .Q(n96) );
  AO22X1 U118 ( .IN1(wr_data[17]), .IN2(n2209), .IN3(\r[1][17] ), .IN4(n2207),
        .Q(n97) );
  AO22X1 U119 ( .IN1(wr_data[18]), .IN2(n2209), .IN3(\r[1][18] ), .IN4(n2207),
        .Q(n98) );
  AO22X1 U120 ( .IN1(wr_data[19]), .IN2(n2209), .IN3(\r[1][19] ), .IN4(n2207),
        .Q(n99) );
  AO22X1 U121 ( .IN1(wr_data[20]), .IN2(n2209), .IN3(\r[1][20] ), .IN4(n2206),
        .Q(n100) );
  AO22X1 U122 ( .IN1(wr_data[21]), .IN2(n2209), .IN3(\r[1][21] ), .IN4(n2206),
        .Q(n101) );
  AO22X1 U123 ( .IN1(wr_data[22]), .IN2(n2209), .IN3(\r[1][22] ), .IN4(n2206),
        .Q(n102) );
  AO22X1 U124 ( .IN1(wr_data[23]), .IN2(n2210), .IN3(\r[1][23] ), .IN4(n2206),
        .Q(n103) );
  AO22X1 U125 ( .IN1(wr_data[24]), .IN2(n2210), .IN3(\r[1][24] ), .IN4(n2206),
        .Q(n104) );
  AO22X1 U126 ( .IN1(wr_data[25]), .IN2(n2210), .IN3(\r[1][25] ), .IN4(n2206),
        .Q(n105) );
  AO22X1 U127 ( .IN1(wr_data[26]), .IN2(n2210), .IN3(\r[1][26] ), .IN4(n2206),
        .Q(n106) );
  AO22X1 U128 ( .IN1(wr_data[27]), .IN2(n2210), .IN3(\r[1][27] ), .IN4(n2206),
        .Q(n107) );
  AO22X1 U129 ( .IN1(wr_data[28]), .IN2(n2210), .IN3(\r[1][28] ), .IN4(n2206),
        .Q(n108) );
  AO22X1 U130 ( .IN1(wr_data[29]), .IN2(n2210), .IN3(\r[1][29] ), .IN4(n2206),
        .Q(n109) );
  AO22X1 U131 ( .IN1(wr_data[30]), .IN2(n2210), .IN3(\r[1][30] ), .IN4(n2206),
        .Q(n110) );
  AO22X1 U132 ( .IN1(wr_data[31]), .IN2(n2210), .IN3(\r[1][31] ), .IN4(n2206),
        .Q(n111) );
  AO22X1 U133 ( .IN1(n2203), .IN2(wr_data[0]), .IN3(\r[2][0] ), .IN4(n40), .Q(
        n112) );
  AO22X1 U134 ( .IN1(n2203), .IN2(wr_data[1]), .IN3(\r[2][1] ), .IN4(n40), .Q(
        n113) );
  AO22X1 U135 ( .IN1(n2203), .IN2(wr_data[2]), .IN3(\r[2][2] ), .IN4(n40), .Q(
        n114) );
  AO22X1 U136 ( .IN1(n2203), .IN2(wr_data[3]), .IN3(\r[2][3] ), .IN4(n40), .Q(
        n115) );
  AO22X1 U137 ( .IN1(n2203), .IN2(wr_data[4]), .IN3(\r[2][4] ), .IN4(n40), .Q(
        n116) );
  AO22X1 U138 ( .IN1(n2203), .IN2(wr_data[5]), .IN3(\r[2][5] ), .IN4(n40), .Q(
        n117) );
  AO22X1 U139 ( .IN1(n2203), .IN2(wr_data[6]), .IN3(\r[2][6] ), .IN4(n40), .Q(
        n118) );
  AO22X1 U140 ( .IN1(n2203), .IN2(wr_data[7]), .IN3(\r[2][7] ), .IN4(n40), .Q(
        n119) );
  AO22X1 U141 ( .IN1(n2203), .IN2(wr_data[8]), .IN3(\r[2][8] ), .IN4(n2202),
        .Q(n120) );
  AO22X1 U142 ( .IN1(n2203), .IN2(wr_data[9]), .IN3(\r[2][9] ), .IN4(n2202),
        .Q(n121) );
  AO22X1 U143 ( .IN1(n2204), .IN2(wr_data[10]), .IN3(\r[2][10] ), .IN4(n2202),
        .Q(n122) );
  AO22X1 U144 ( .IN1(n2204), .IN2(wr_data[11]), .IN3(\r[2][11] ), .IN4(n2202),
        .Q(n123) );
  AO22X1 U145 ( .IN1(n2204), .IN2(wr_data[12]), .IN3(\r[2][12] ), .IN4(n2202),
        .Q(n124) );
  AO22X1 U146 ( .IN1(n2204), .IN2(wr_data[13]), .IN3(\r[2][13] ), .IN4(n2202),
        .Q(n125) );
  AO22X1 U147 ( .IN1(n2204), .IN2(wr_data[14]), .IN3(\r[2][14] ), .IN4(n2202),
        .Q(n126) );
  AO22X1 U148 ( .IN1(n2204), .IN2(wr_data[15]), .IN3(\r[2][15] ), .IN4(n2202),
        .Q(n127) );
  AO22X1 U149 ( .IN1(n2204), .IN2(wr_data[16]), .IN3(\r[2][16] ), .IN4(n2202),
        .Q(n128) );
  AO22X1 U150 ( .IN1(n2204), .IN2(wr_data[17]), .IN3(\r[2][17] ), .IN4(n2202),
        .Q(n129) );
  AO22X1 U151 ( .IN1(n2204), .IN2(wr_data[18]), .IN3(\r[2][18] ), .IN4(n2202),
        .Q(n130) );
  AO22X1 U152 ( .IN1(n2204), .IN2(wr_data[19]), .IN3(\r[2][19] ), .IN4(n2202),
        .Q(n131) );
  AO22X1 U153 ( .IN1(n2204), .IN2(wr_data[20]), .IN3(\r[2][20] ), .IN4(n2201),
        .Q(n132) );
  AO22X1 U154 ( .IN1(n2204), .IN2(wr_data[21]), .IN3(\r[2][21] ), .IN4(n2201),
        .Q(n133) );
  AO22X1 U155 ( .IN1(n2204), .IN2(wr_data[22]), .IN3(\r[2][22] ), .IN4(n2201),
        .Q(n134) );
  AO22X1 U156 ( .IN1(n2205), .IN2(wr_data[23]), .IN3(\r[2][23] ), .IN4(n2201),
        .Q(n135) );
  AO22X1 U157 ( .IN1(n2205), .IN2(wr_data[24]), .IN3(\r[2][24] ), .IN4(n2201),
        .Q(n136) );
  AO22X1 U158 ( .IN1(n2205), .IN2(wr_data[25]), .IN3(\r[2][25] ), .IN4(n2201),
        .Q(n137) );
  AO22X1 U159 ( .IN1(n2205), .IN2(wr_data[26]), .IN3(\r[2][26] ), .IN4(n2201),
        .Q(n138) );
  AO22X1 U160 ( .IN1(n2205), .IN2(wr_data[27]), .IN3(\r[2][27] ), .IN4(n2201),
        .Q(n139) );
  AO22X1 U161 ( .IN1(n2205), .IN2(wr_data[28]), .IN3(\r[2][28] ), .IN4(n2201),
        .Q(n140) );
  AO22X1 U162 ( .IN1(n2205), .IN2(wr_data[29]), .IN3(\r[2][29] ), .IN4(n2201),
        .Q(n141) );
  AO22X1 U163 ( .IN1(n2205), .IN2(wr_data[30]), .IN3(\r[2][30] ), .IN4(n2201),
        .Q(n142) );
  AO22X1 U164 ( .IN1(n2205), .IN2(wr_data[31]), .IN3(\r[2][31] ), .IN4(n2201),
        .Q(n143) );
  AO22X1 U165 ( .IN1(n2198), .IN2(wr_data[0]), .IN3(\r[3][0] ), .IN4(n42), .Q(
        n144) );
  AO22X1 U166 ( .IN1(n2198), .IN2(wr_data[1]), .IN3(\r[3][1] ), .IN4(n42), .Q(
        n145) );
  AO22X1 U167 ( .IN1(n2198), .IN2(wr_data[2]), .IN3(\r[3][2] ), .IN4(n42), .Q(
        n146) );
  AO22X1 U168 ( .IN1(n2198), .IN2(wr_data[3]), .IN3(\r[3][3] ), .IN4(n42), .Q(
        n147) );
  AO22X1 U169 ( .IN1(n2198), .IN2(wr_data[4]), .IN3(\r[3][4] ), .IN4(n42), .Q(
        n148) );
  AO22X1 U170 ( .IN1(n2198), .IN2(wr_data[5]), .IN3(\r[3][5] ), .IN4(n42), .Q(
        n149) );
  AO22X1 U171 ( .IN1(n2198), .IN2(wr_data[6]), .IN3(\r[3][6] ), .IN4(n42), .Q(
        n150) );
  AO22X1 U172 ( .IN1(n2198), .IN2(wr_data[7]), .IN3(\r[3][7] ), .IN4(n42), .Q(
        n151) );
  AO22X1 U173 ( .IN1(n2198), .IN2(wr_data[8]), .IN3(\r[3][8] ), .IN4(n2197),
        .Q(n152) );
  AO22X1 U174 ( .IN1(n2198), .IN2(wr_data[9]), .IN3(\r[3][9] ), .IN4(n2197),
        .Q(n153) );
  AO22X1 U175 ( .IN1(n2199), .IN2(wr_data[10]), .IN3(\r[3][10] ), .IN4(n2197),
        .Q(n154) );
  AO22X1 U176 ( .IN1(n2199), .IN2(wr_data[11]), .IN3(\r[3][11] ), .IN4(n2197),
        .Q(n155) );
  AO22X1 U177 ( .IN1(n2199), .IN2(wr_data[12]), .IN3(\r[3][12] ), .IN4(n2197),
        .Q(n156) );
  AO22X1 U178 ( .IN1(n2199), .IN2(wr_data[13]), .IN3(\r[3][13] ), .IN4(n2197),
        .Q(n157) );
  AO22X1 U179 ( .IN1(n2199), .IN2(wr_data[14]), .IN3(\r[3][14] ), .IN4(n2197),
        .Q(n158) );
  AO22X1 U180 ( .IN1(n2199), .IN2(wr_data[15]), .IN3(\r[3][15] ), .IN4(n2197),
        .Q(n159) );
  AO22X1 U181 ( .IN1(n2199), .IN2(wr_data[16]), .IN3(\r[3][16] ), .IN4(n2197),
        .Q(n160) );
  AO22X1 U182 ( .IN1(n2199), .IN2(wr_data[17]), .IN3(\r[3][17] ), .IN4(n2197),
        .Q(n161) );
  AO22X1 U183 ( .IN1(n2199), .IN2(wr_data[18]), .IN3(\r[3][18] ), .IN4(n2197),
        .Q(n162) );
  AO22X1 U184 ( .IN1(n2199), .IN2(wr_data[19]), .IN3(\r[3][19] ), .IN4(n2197),
        .Q(n163) );
  AO22X1 U185 ( .IN1(n2199), .IN2(wr_data[20]), .IN3(\r[3][20] ), .IN4(n2196),
        .Q(n164) );
  AO22X1 U186 ( .IN1(n2199), .IN2(wr_data[21]), .IN3(\r[3][21] ), .IN4(n2196),
        .Q(n165) );
  AO22X1 U187 ( .IN1(n2199), .IN2(wr_data[22]), .IN3(\r[3][22] ), .IN4(n2196),
        .Q(n166) );
  AO22X1 U188 ( .IN1(n2200), .IN2(wr_data[23]), .IN3(\r[3][23] ), .IN4(n2196),
        .Q(n167) );
  AO22X1 U189 ( .IN1(n2200), .IN2(wr_data[24]), .IN3(\r[3][24] ), .IN4(n2196),
        .Q(n168) );
  AO22X1 U190 ( .IN1(n2200), .IN2(wr_data[25]), .IN3(\r[3][25] ), .IN4(n2196),
        .Q(n169) );
  AO22X1 U191 ( .IN1(n2200), .IN2(wr_data[26]), .IN3(\r[3][26] ), .IN4(n2196),
        .Q(n170) );
  AO22X1 U192 ( .IN1(n2200), .IN2(wr_data[27]), .IN3(\r[3][27] ), .IN4(n2196),
        .Q(n171) );
  AO22X1 U193 ( .IN1(n2200), .IN2(wr_data[28]), .IN3(\r[3][28] ), .IN4(n2196),
        .Q(n172) );
  AO22X1 U194 ( .IN1(n2200), .IN2(wr_data[29]), .IN3(\r[3][29] ), .IN4(n2196),
        .Q(n173) );
  AO22X1 U195 ( .IN1(n2200), .IN2(wr_data[30]), .IN3(\r[3][30] ), .IN4(n2196),
        .Q(n174) );
  AO22X1 U196 ( .IN1(n2200), .IN2(wr_data[31]), .IN3(\r[3][31] ), .IN4(n2196),
        .Q(n175) );
  AO22X1 U197 ( .IN1(n2193), .IN2(wr_data[0]), .IN3(\r[4][0] ), .IN4(n44), .Q(
        n176) );
  AO22X1 U198 ( .IN1(n2193), .IN2(wr_data[1]), .IN3(\r[4][1] ), .IN4(n44), .Q(
        n177) );
  AO22X1 U199 ( .IN1(n2193), .IN2(wr_data[2]), .IN3(\r[4][2] ), .IN4(n44), .Q(
        n178) );
  AO22X1 U200 ( .IN1(n2193), .IN2(wr_data[3]), .IN3(\r[4][3] ), .IN4(n44), .Q(
        n179) );
  AO22X1 U201 ( .IN1(n2193), .IN2(wr_data[4]), .IN3(\r[4][4] ), .IN4(n44), .Q(
        n180) );
  AO22X1 U202 ( .IN1(n2193), .IN2(wr_data[5]), .IN3(\r[4][5] ), .IN4(n44), .Q(
        n181) );
  AO22X1 U203 ( .IN1(n2193), .IN2(wr_data[6]), .IN3(\r[4][6] ), .IN4(n44), .Q(
        n182) );
  AO22X1 U204 ( .IN1(n2193), .IN2(wr_data[7]), .IN3(\r[4][7] ), .IN4(n44), .Q(
        n183) );
  AO22X1 U205 ( .IN1(n2193), .IN2(wr_data[8]), .IN3(\r[4][8] ), .IN4(n2192),
        .Q(n184) );
  AO22X1 U206 ( .IN1(n2193), .IN2(wr_data[9]), .IN3(\r[4][9] ), .IN4(n2192),
        .Q(n185) );
  AO22X1 U207 ( .IN1(n2194), .IN2(wr_data[10]), .IN3(\r[4][10] ), .IN4(n2192),
        .Q(n186) );
  AO22X1 U208 ( .IN1(n2194), .IN2(wr_data[11]), .IN3(\r[4][11] ), .IN4(n2192),
        .Q(n187) );
  AO22X1 U209 ( .IN1(n2194), .IN2(wr_data[12]), .IN3(\r[4][12] ), .IN4(n2192),
        .Q(n188) );
  AO22X1 U210 ( .IN1(n2194), .IN2(wr_data[13]), .IN3(\r[4][13] ), .IN4(n2192),
        .Q(n189) );
  AO22X1 U211 ( .IN1(n2194), .IN2(wr_data[14]), .IN3(\r[4][14] ), .IN4(n2192),
        .Q(n190) );
  AO22X1 U212 ( .IN1(n2194), .IN2(wr_data[15]), .IN3(\r[4][15] ), .IN4(n2192),
        .Q(n191) );
  AO22X1 U213 ( .IN1(n2194), .IN2(wr_data[16]), .IN3(\r[4][16] ), .IN4(n2192),
        .Q(n192) );
  AO22X1 U214 ( .IN1(n2194), .IN2(wr_data[17]), .IN3(\r[4][17] ), .IN4(n2192),
        .Q(n193) );
  AO22X1 U215 ( .IN1(n2194), .IN2(wr_data[18]), .IN3(\r[4][18] ), .IN4(n2192),
        .Q(n194) );
  AO22X1 U216 ( .IN1(n2194), .IN2(wr_data[19]), .IN3(\r[4][19] ), .IN4(n2192),
        .Q(n195) );
  AO22X1 U217 ( .IN1(n2194), .IN2(wr_data[20]), .IN3(\r[4][20] ), .IN4(n2191),
        .Q(n196) );
  AO22X1 U218 ( .IN1(n2194), .IN2(wr_data[21]), .IN3(\r[4][21] ), .IN4(n2191),
        .Q(n197) );
  AO22X1 U219 ( .IN1(n2194), .IN2(wr_data[22]), .IN3(\r[4][22] ), .IN4(n2191),
        .Q(n198) );
  AO22X1 U220 ( .IN1(n2195), .IN2(wr_data[23]), .IN3(\r[4][23] ), .IN4(n2191),
        .Q(n199) );
  AO22X1 U221 ( .IN1(n2195), .IN2(wr_data[24]), .IN3(\r[4][24] ), .IN4(n2191),
        .Q(n200) );
  AO22X1 U222 ( .IN1(n2195), .IN2(wr_data[25]), .IN3(\r[4][25] ), .IN4(n2191),
        .Q(n201) );
  AO22X1 U223 ( .IN1(n2195), .IN2(wr_data[26]), .IN3(\r[4][26] ), .IN4(n2191),
        .Q(n202) );
  AO22X1 U224 ( .IN1(n2195), .IN2(wr_data[27]), .IN3(\r[4][27] ), .IN4(n2191),
        .Q(n203) );
  AO22X1 U225 ( .IN1(n2195), .IN2(wr_data[28]), .IN3(\r[4][28] ), .IN4(n2191),
        .Q(n204) );
  AO22X1 U226 ( .IN1(n2195), .IN2(wr_data[29]), .IN3(\r[4][29] ), .IN4(n2191),
        .Q(n205) );
  AO22X1 U227 ( .IN1(n2195), .IN2(wr_data[30]), .IN3(\r[4][30] ), .IN4(n2191),
        .Q(n206) );
  AO22X1 U228 ( .IN1(n2195), .IN2(wr_data[31]), .IN3(\r[4][31] ), .IN4(n2191),
        .Q(n207) );
  AO22X1 U229 ( .IN1(n2188), .IN2(wr_data[0]), .IN3(\r[5][0] ), .IN4(n46), .Q(
        n208) );
  AO22X1 U230 ( .IN1(n2188), .IN2(wr_data[1]), .IN3(\r[5][1] ), .IN4(n46), .Q(
        n209) );
  AO22X1 U231 ( .IN1(n2188), .IN2(wr_data[2]), .IN3(\r[5][2] ), .IN4(n46), .Q(
        n210) );
  AO22X1 U232 ( .IN1(n2188), .IN2(wr_data[3]), .IN3(\r[5][3] ), .IN4(n46), .Q(
        n211) );
  AO22X1 U233 ( .IN1(n2188), .IN2(wr_data[4]), .IN3(\r[5][4] ), .IN4(n46), .Q(
        n212) );
  AO22X1 U234 ( .IN1(n2188), .IN2(wr_data[5]), .IN3(\r[5][5] ), .IN4(n46), .Q(
        n213) );
  AO22X1 U235 ( .IN1(n2188), .IN2(wr_data[6]), .IN3(\r[5][6] ), .IN4(n46), .Q(
        n214) );
  AO22X1 U236 ( .IN1(n2188), .IN2(wr_data[7]), .IN3(\r[5][7] ), .IN4(n46), .Q(
        n215) );
  AO22X1 U237 ( .IN1(n2188), .IN2(wr_data[8]), .IN3(\r[5][8] ), .IN4(n2187),
        .Q(n216) );
  AO22X1 U238 ( .IN1(n2188), .IN2(wr_data[9]), .IN3(\r[5][9] ), .IN4(n2187),
        .Q(n217) );
  AO22X1 U239 ( .IN1(n2189), .IN2(wr_data[10]), .IN3(\r[5][10] ), .IN4(n2187),
        .Q(n218) );
  AO22X1 U240 ( .IN1(n2189), .IN2(wr_data[11]), .IN3(\r[5][11] ), .IN4(n2187),
        .Q(n219) );
  AO22X1 U241 ( .IN1(n2189), .IN2(wr_data[12]), .IN3(\r[5][12] ), .IN4(n2187),
        .Q(n220) );
  AO22X1 U242 ( .IN1(n2189), .IN2(wr_data[13]), .IN3(\r[5][13] ), .IN4(n2187),
        .Q(n221) );
  AO22X1 U243 ( .IN1(n2189), .IN2(wr_data[14]), .IN3(\r[5][14] ), .IN4(n2187),
        .Q(n222) );
  AO22X1 U244 ( .IN1(n2189), .IN2(wr_data[15]), .IN3(\r[5][15] ), .IN4(n2187),
        .Q(n223) );
  AO22X1 U245 ( .IN1(n2189), .IN2(wr_data[16]), .IN3(\r[5][16] ), .IN4(n2187),
        .Q(n224) );
  AO22X1 U246 ( .IN1(n2189), .IN2(wr_data[17]), .IN3(\r[5][17] ), .IN4(n2187),
        .Q(n225) );
  AO22X1 U247 ( .IN1(n2189), .IN2(wr_data[18]), .IN3(\r[5][18] ), .IN4(n2187),
        .Q(n226) );
  AO22X1 U248 ( .IN1(n2189), .IN2(wr_data[19]), .IN3(\r[5][19] ), .IN4(n2187),
        .Q(n227) );
  AO22X1 U249 ( .IN1(n2189), .IN2(wr_data[20]), .IN3(\r[5][20] ), .IN4(n2186),
        .Q(n228) );
  AO22X1 U250 ( .IN1(n2189), .IN2(wr_data[21]), .IN3(\r[5][21] ), .IN4(n2186),
        .Q(n229) );
  AO22X1 U251 ( .IN1(n2189), .IN2(wr_data[22]), .IN3(\r[5][22] ), .IN4(n2186),
        .Q(n230) );
  AO22X1 U252 ( .IN1(n2190), .IN2(wr_data[23]), .IN3(\r[5][23] ), .IN4(n2186),
        .Q(n231) );
  AO22X1 U253 ( .IN1(n2190), .IN2(wr_data[24]), .IN3(\r[5][24] ), .IN4(n2186),
        .Q(n232) );
  AO22X1 U254 ( .IN1(n2190), .IN2(wr_data[25]), .IN3(\r[5][25] ), .IN4(n2186),
        .Q(n233) );
  AO22X1 U255 ( .IN1(n2190), .IN2(wr_data[26]), .IN3(\r[5][26] ), .IN4(n2186),
        .Q(n234) );
  AO22X1 U256 ( .IN1(n2190), .IN2(wr_data[27]), .IN3(\r[5][27] ), .IN4(n2186),
        .Q(n235) );
  AO22X1 U257 ( .IN1(n2190), .IN2(wr_data[28]), .IN3(\r[5][28] ), .IN4(n2186),
        .Q(n236) );
  AO22X1 U258 ( .IN1(n2190), .IN2(wr_data[29]), .IN3(\r[5][29] ), .IN4(n2186),
        .Q(n237) );
  AO22X1 U259 ( .IN1(n2190), .IN2(wr_data[30]), .IN3(\r[5][30] ), .IN4(n2186),
        .Q(n238) );
  AO22X1 U260 ( .IN1(n2190), .IN2(wr_data[31]), .IN3(\r[5][31] ), .IN4(n2186),
        .Q(n239) );
  AO22X1 U261 ( .IN1(n2183), .IN2(wr_data[0]), .IN3(\r[6][0] ), .IN4(n48), .Q(
        n240) );
  AO22X1 U262 ( .IN1(n2183), .IN2(wr_data[1]), .IN3(\r[6][1] ), .IN4(n48), .Q(
        n241) );
  AO22X1 U263 ( .IN1(n2183), .IN2(wr_data[2]), .IN3(\r[6][2] ), .IN4(n48), .Q(
        n242) );
  AO22X1 U264 ( .IN1(n2183), .IN2(wr_data[3]), .IN3(\r[6][3] ), .IN4(n48), .Q(
        n243) );
  AO22X1 U265 ( .IN1(n2183), .IN2(wr_data[4]), .IN3(\r[6][4] ), .IN4(n48), .Q(
        n244) );
  AO22X1 U266 ( .IN1(n2183), .IN2(wr_data[5]), .IN3(\r[6][5] ), .IN4(n48), .Q(
        n245) );
  AO22X1 U267 ( .IN1(n2183), .IN2(wr_data[6]), .IN3(\r[6][6] ), .IN4(n48), .Q(
        n246) );
  AO22X1 U268 ( .IN1(n2183), .IN2(wr_data[7]), .IN3(\r[6][7] ), .IN4(n48), .Q(
        n247) );
  AO22X1 U269 ( .IN1(n2183), .IN2(wr_data[8]), .IN3(\r[6][8] ), .IN4(n2182),
        .Q(n248) );
  AO22X1 U270 ( .IN1(n2183), .IN2(wr_data[9]), .IN3(\r[6][9] ), .IN4(n2182),
        .Q(n249) );
  AO22X1 U271 ( .IN1(n2184), .IN2(wr_data[10]), .IN3(\r[6][10] ), .IN4(n2182),
        .Q(n250) );
  AO22X1 U272 ( .IN1(n2184), .IN2(wr_data[11]), .IN3(\r[6][11] ), .IN4(n2182),
        .Q(n251) );
  AO22X1 U273 ( .IN1(n2184), .IN2(wr_data[12]), .IN3(\r[6][12] ), .IN4(n2182),
        .Q(n252) );
  AO22X1 U274 ( .IN1(n2184), .IN2(wr_data[13]), .IN3(\r[6][13] ), .IN4(n2182),
        .Q(n253) );
  AO22X1 U275 ( .IN1(n2184), .IN2(wr_data[14]), .IN3(\r[6][14] ), .IN4(n2182),
        .Q(n254) );
  AO22X1 U276 ( .IN1(n2184), .IN2(wr_data[15]), .IN3(\r[6][15] ), .IN4(n2182),
        .Q(n255) );
  AO22X1 U277 ( .IN1(n2184), .IN2(wr_data[16]), .IN3(\r[6][16] ), .IN4(n2182),
        .Q(n256) );
  AO22X1 U278 ( .IN1(n2184), .IN2(wr_data[17]), .IN3(\r[6][17] ), .IN4(n2182),
        .Q(n257) );
  AO22X1 U279 ( .IN1(n2184), .IN2(wr_data[18]), .IN3(\r[6][18] ), .IN4(n2182),
        .Q(n258) );
  AO22X1 U280 ( .IN1(n2184), .IN2(wr_data[19]), .IN3(\r[6][19] ), .IN4(n2182),
        .Q(n259) );
  AO22X1 U281 ( .IN1(n2184), .IN2(wr_data[20]), .IN3(\r[6][20] ), .IN4(n2181),
        .Q(n260) );
  AO22X1 U282 ( .IN1(n2184), .IN2(wr_data[21]), .IN3(\r[6][21] ), .IN4(n2181),
        .Q(n261) );
  AO22X1 U283 ( .IN1(n2184), .IN2(wr_data[22]), .IN3(\r[6][22] ), .IN4(n2181),
        .Q(n262) );
  AO22X1 U284 ( .IN1(n2185), .IN2(wr_data[23]), .IN3(\r[6][23] ), .IN4(n2181),
        .Q(n263) );
  AO22X1 U285 ( .IN1(n2185), .IN2(wr_data[24]), .IN3(\r[6][24] ), .IN4(n2181),
        .Q(n264) );
  AO22X1 U286 ( .IN1(n2185), .IN2(wr_data[25]), .IN3(\r[6][25] ), .IN4(n2181),
        .Q(n265) );
  AO22X1 U287 ( .IN1(n2185), .IN2(wr_data[26]), .IN3(\r[6][26] ), .IN4(n2181),
        .Q(n266) );
  AO22X1 U288 ( .IN1(n2185), .IN2(wr_data[27]), .IN3(\r[6][27] ), .IN4(n2181),
        .Q(n267) );
  AO22X1 U289 ( .IN1(n2185), .IN2(wr_data[28]), .IN3(\r[6][28] ), .IN4(n2181),
        .Q(n268) );
  AO22X1 U290 ( .IN1(n2185), .IN2(wr_data[29]), .IN3(\r[6][29] ), .IN4(n2181),
        .Q(n269) );
  AO22X1 U291 ( .IN1(n2185), .IN2(wr_data[30]), .IN3(\r[6][30] ), .IN4(n2181),
        .Q(n270) );
  AO22X1 U292 ( .IN1(n2185), .IN2(wr_data[31]), .IN3(\r[6][31] ), .IN4(n2181),
        .Q(n271) );
  AO22X1 U293 ( .IN1(n2178), .IN2(wr_data[0]), .IN3(\r[7][0] ), .IN4(n50), .Q(
        n272) );
  AO22X1 U294 ( .IN1(n2178), .IN2(wr_data[1]), .IN3(\r[7][1] ), .IN4(n50), .Q(
        n273) );
  AO22X1 U295 ( .IN1(n2178), .IN2(wr_data[2]), .IN3(\r[7][2] ), .IN4(n50), .Q(
        n274) );
  AO22X1 U296 ( .IN1(n2178), .IN2(wr_data[3]), .IN3(\r[7][3] ), .IN4(n50), .Q(
        n275) );
  AO22X1 U297 ( .IN1(n2178), .IN2(wr_data[4]), .IN3(\r[7][4] ), .IN4(n50), .Q(
        n276) );
  AO22X1 U298 ( .IN1(n2178), .IN2(wr_data[5]), .IN3(\r[7][5] ), .IN4(n50), .Q(
        n277) );
  AO22X1 U299 ( .IN1(n2178), .IN2(wr_data[6]), .IN3(\r[7][6] ), .IN4(n50), .Q(
        n278) );
  AO22X1 U300 ( .IN1(n2178), .IN2(wr_data[7]), .IN3(\r[7][7] ), .IN4(n50), .Q(
        n279) );
  AO22X1 U301 ( .IN1(n2178), .IN2(wr_data[8]), .IN3(\r[7][8] ), .IN4(n2177),
        .Q(n280) );
  AO22X1 U302 ( .IN1(n2178), .IN2(wr_data[9]), .IN3(\r[7][9] ), .IN4(n2177),
        .Q(n281) );
  AO22X1 U303 ( .IN1(n2179), .IN2(wr_data[10]), .IN3(\r[7][10] ), .IN4(n2177),
        .Q(n282) );
  AO22X1 U304 ( .IN1(n2179), .IN2(wr_data[11]), .IN3(\r[7][11] ), .IN4(n2177),
        .Q(n283) );
  AO22X1 U305 ( .IN1(n2179), .IN2(wr_data[12]), .IN3(\r[7][12] ), .IN4(n2177),
        .Q(n284) );
  AO22X1 U306 ( .IN1(n2179), .IN2(wr_data[13]), .IN3(\r[7][13] ), .IN4(n2177),
        .Q(n285) );
  AO22X1 U307 ( .IN1(n2179), .IN2(wr_data[14]), .IN3(\r[7][14] ), .IN4(n2177),
        .Q(n286) );
  AO22X1 U308 ( .IN1(n2179), .IN2(wr_data[15]), .IN3(\r[7][15] ), .IN4(n2177),
        .Q(n287) );
  AO22X1 U309 ( .IN1(n2179), .IN2(wr_data[16]), .IN3(\r[7][16] ), .IN4(n2177),
        .Q(n288) );
  AO22X1 U310 ( .IN1(n2179), .IN2(wr_data[17]), .IN3(\r[7][17] ), .IN4(n2177),
        .Q(n289) );
  AO22X1 U311 ( .IN1(n2179), .IN2(wr_data[18]), .IN3(\r[7][18] ), .IN4(n2177),
        .Q(n290) );
  AO22X1 U312 ( .IN1(n2179), .IN2(wr_data[19]), .IN3(\r[7][19] ), .IN4(n2177),
        .Q(n291) );
  AO22X1 U313 ( .IN1(n2179), .IN2(wr_data[20]), .IN3(\r[7][20] ), .IN4(n2176),
        .Q(n292) );
  AO22X1 U314 ( .IN1(n2179), .IN2(wr_data[21]), .IN3(\r[7][21] ), .IN4(n2176),
        .Q(n293) );
  AO22X1 U315 ( .IN1(n2179), .IN2(wr_data[22]), .IN3(\r[7][22] ), .IN4(n2176),
        .Q(n294) );
  AO22X1 U316 ( .IN1(n2180), .IN2(wr_data[23]), .IN3(\r[7][23] ), .IN4(n2176),
        .Q(n295) );
  AO22X1 U317 ( .IN1(n2180), .IN2(wr_data[24]), .IN3(\r[7][24] ), .IN4(n2176),
        .Q(n296) );
  AO22X1 U318 ( .IN1(n2180), .IN2(wr_data[25]), .IN3(\r[7][25] ), .IN4(n2176),
        .Q(n297) );
  AO22X1 U319 ( .IN1(n2180), .IN2(wr_data[26]), .IN3(\r[7][26] ), .IN4(n2176),
        .Q(n298) );
  AO22X1 U320 ( .IN1(n2180), .IN2(wr_data[27]), .IN3(\r[7][27] ), .IN4(n2176),
        .Q(n299) );
  AO22X1 U321 ( .IN1(n2180), .IN2(wr_data[28]), .IN3(\r[7][28] ), .IN4(n2176),
        .Q(n300) );
  AO22X1 U322 ( .IN1(n2180), .IN2(wr_data[29]), .IN3(\r[7][29] ), .IN4(n2176),
        .Q(n301) );
  AO22X1 U323 ( .IN1(n2180), .IN2(wr_data[30]), .IN3(\r[7][30] ), .IN4(n2176),
        .Q(n302) );
  AO22X1 U324 ( .IN1(n2180), .IN2(wr_data[31]), .IN3(\r[7][31] ), .IN4(n2176),
        .Q(n303) );
  AND3X1 U325 ( .IN1(n2300), .IN2(n2299), .IN3(wr_en), .Q(n39) );
  AO22X1 U326 ( .IN1(n2173), .IN2(wr_data[0]), .IN3(\r[8][0] ), .IN4(n52), .Q(
        n304) );
  AO22X1 U327 ( .IN1(n2173), .IN2(wr_data[1]), .IN3(\r[8][1] ), .IN4(n52), .Q(
        n305) );
  AO22X1 U328 ( .IN1(n2173), .IN2(wr_data[2]), .IN3(\r[8][2] ), .IN4(n52), .Q(
        n306) );
  AO22X1 U329 ( .IN1(n2173), .IN2(wr_data[3]), .IN3(\r[8][3] ), .IN4(n52), .Q(
        n307) );
  AO22X1 U330 ( .IN1(n2173), .IN2(wr_data[4]), .IN3(\r[8][4] ), .IN4(n52), .Q(
        n308) );
  AO22X1 U331 ( .IN1(n2173), .IN2(wr_data[5]), .IN3(\r[8][5] ), .IN4(n52), .Q(
        n309) );
  AO22X1 U332 ( .IN1(n2173), .IN2(wr_data[6]), .IN3(\r[8][6] ), .IN4(n52), .Q(
        n310) );
  AO22X1 U333 ( .IN1(n2173), .IN2(wr_data[7]), .IN3(\r[8][7] ), .IN4(n52), .Q(
        n311) );
  AO22X1 U334 ( .IN1(n2173), .IN2(wr_data[8]), .IN3(\r[8][8] ), .IN4(n2172),
        .Q(n312) );
  AO22X1 U335 ( .IN1(n2173), .IN2(wr_data[9]), .IN3(\r[8][9] ), .IN4(n2172),
        .Q(n313) );
  AO22X1 U336 ( .IN1(n2174), .IN2(wr_data[10]), .IN3(\r[8][10] ), .IN4(n2172),
        .Q(n314) );
  AO22X1 U337 ( .IN1(n2174), .IN2(wr_data[11]), .IN3(\r[8][11] ), .IN4(n2172),
        .Q(n315) );
  AO22X1 U338 ( .IN1(n2174), .IN2(wr_data[12]), .IN3(\r[8][12] ), .IN4(n2172),
        .Q(n316) );
  AO22X1 U339 ( .IN1(n2174), .IN2(wr_data[13]), .IN3(\r[8][13] ), .IN4(n2172),
        .Q(n317) );
  AO22X1 U340 ( .IN1(n2174), .IN2(wr_data[14]), .IN3(\r[8][14] ), .IN4(n2172),
        .Q(n318) );
  AO22X1 U341 ( .IN1(n2174), .IN2(wr_data[15]), .IN3(\r[8][15] ), .IN4(n2172),
        .Q(n319) );
  AO22X1 U342 ( .IN1(n2174), .IN2(wr_data[16]), .IN3(\r[8][16] ), .IN4(n2172),
        .Q(n320) );
  AO22X1 U343 ( .IN1(n2174), .IN2(wr_data[17]), .IN3(\r[8][17] ), .IN4(n2172),
        .Q(n321) );
  AO22X1 U344 ( .IN1(n2174), .IN2(wr_data[18]), .IN3(\r[8][18] ), .IN4(n2172),
        .Q(n322) );
  AO22X1 U345 ( .IN1(n2174), .IN2(wr_data[19]), .IN3(\r[8][19] ), .IN4(n2172),
        .Q(n323) );
  AO22X1 U346 ( .IN1(n2174), .IN2(wr_data[20]), .IN3(\r[8][20] ), .IN4(n2171),
        .Q(n324) );
  AO22X1 U347 ( .IN1(n2174), .IN2(wr_data[21]), .IN3(\r[8][21] ), .IN4(n2171),
        .Q(n325) );
  AO22X1 U348 ( .IN1(n2174), .IN2(wr_data[22]), .IN3(\r[8][22] ), .IN4(n2171),
        .Q(n326) );
  AO22X1 U349 ( .IN1(n2175), .IN2(wr_data[23]), .IN3(\r[8][23] ), .IN4(n2171),
        .Q(n327) );
  AO22X1 U350 ( .IN1(n2175), .IN2(wr_data[24]), .IN3(\r[8][24] ), .IN4(n2171),
        .Q(n328) );
  AO22X1 U351 ( .IN1(n2175), .IN2(wr_data[25]), .IN3(\r[8][25] ), .IN4(n2171),
        .Q(n329) );
  AO22X1 U352 ( .IN1(n2175), .IN2(wr_data[26]), .IN3(\r[8][26] ), .IN4(n2171),
        .Q(n330) );
  AO22X1 U353 ( .IN1(n2175), .IN2(wr_data[27]), .IN3(\r[8][27] ), .IN4(n2171),
        .Q(n331) );
  AO22X1 U354 ( .IN1(n2175), .IN2(wr_data[28]), .IN3(\r[8][28] ), .IN4(n2171),
        .Q(n332) );
  AO22X1 U355 ( .IN1(n2175), .IN2(wr_data[29]), .IN3(\r[8][29] ), .IN4(n2171),
        .Q(n333) );
  AO22X1 U356 ( .IN1(n2175), .IN2(wr_data[30]), .IN3(\r[8][30] ), .IN4(n2171),
        .Q(n334) );
  AO22X1 U357 ( .IN1(n2175), .IN2(wr_data[31]), .IN3(\r[8][31] ), .IN4(n2171),
        .Q(n335) );
  AO22X1 U358 ( .IN1(n2168), .IN2(wr_data[0]), .IN3(\r[9][0] ), .IN4(n55), .Q(
        n336) );
  AO22X1 U359 ( .IN1(n2168), .IN2(wr_data[1]), .IN3(\r[9][1] ), .IN4(n55), .Q(
        n337) );
  AO22X1 U360 ( .IN1(n2168), .IN2(wr_data[2]), .IN3(\r[9][2] ), .IN4(n55), .Q(
        n338) );
  AO22X1 U361 ( .IN1(n2168), .IN2(wr_data[3]), .IN3(\r[9][3] ), .IN4(n55), .Q(
        n339) );
  AO22X1 U362 ( .IN1(n2168), .IN2(wr_data[4]), .IN3(\r[9][4] ), .IN4(n55), .Q(
        n340) );
  AO22X1 U363 ( .IN1(n2168), .IN2(wr_data[5]), .IN3(\r[9][5] ), .IN4(n55), .Q(
        n341) );
  AO22X1 U364 ( .IN1(n2168), .IN2(wr_data[6]), .IN3(\r[9][6] ), .IN4(n55), .Q(
        n342) );
  AO22X1 U365 ( .IN1(n2168), .IN2(wr_data[7]), .IN3(\r[9][7] ), .IN4(n55), .Q(
        n343) );
  AO22X1 U366 ( .IN1(n2168), .IN2(wr_data[8]), .IN3(\r[9][8] ), .IN4(n2167),
        .Q(n344) );
  AO22X1 U367 ( .IN1(n2168), .IN2(wr_data[9]), .IN3(\r[9][9] ), .IN4(n2167),
        .Q(n345) );
  AO22X1 U368 ( .IN1(n2169), .IN2(wr_data[10]), .IN3(\r[9][10] ), .IN4(n2167),
        .Q(n346) );
  AO22X1 U369 ( .IN1(n2169), .IN2(wr_data[11]), .IN3(\r[9][11] ), .IN4(n2167),
        .Q(n347) );
  AO22X1 U370 ( .IN1(n2169), .IN2(wr_data[12]), .IN3(\r[9][12] ), .IN4(n2167),
        .Q(n348) );
  AO22X1 U371 ( .IN1(n2169), .IN2(wr_data[13]), .IN3(\r[9][13] ), .IN4(n2167),
        .Q(n349) );
  AO22X1 U372 ( .IN1(n2169), .IN2(wr_data[14]), .IN3(\r[9][14] ), .IN4(n2167),
        .Q(n350) );
  AO22X1 U373 ( .IN1(n2169), .IN2(wr_data[15]), .IN3(\r[9][15] ), .IN4(n2167),
        .Q(n351) );
  AO22X1 U374 ( .IN1(n2169), .IN2(wr_data[16]), .IN3(\r[9][16] ), .IN4(n2167),
        .Q(n352) );
  AO22X1 U375 ( .IN1(n2169), .IN2(wr_data[17]), .IN3(\r[9][17] ), .IN4(n2167),
        .Q(n353) );
  AO22X1 U376 ( .IN1(n2169), .IN2(wr_data[18]), .IN3(\r[9][18] ), .IN4(n2167),
        .Q(n354) );
  AO22X1 U377 ( .IN1(n2169), .IN2(wr_data[19]), .IN3(\r[9][19] ), .IN4(n2167),
        .Q(n355) );
  AO22X1 U378 ( .IN1(n2169), .IN2(wr_data[20]), .IN3(\r[9][20] ), .IN4(n2166),
        .Q(n356) );
  AO22X1 U379 ( .IN1(n2169), .IN2(wr_data[21]), .IN3(\r[9][21] ), .IN4(n2166),
        .Q(n357) );
  AO22X1 U380 ( .IN1(n2169), .IN2(wr_data[22]), .IN3(\r[9][22] ), .IN4(n2166),
        .Q(n358) );
  AO22X1 U381 ( .IN1(n2170), .IN2(wr_data[23]), .IN3(\r[9][23] ), .IN4(n2166),
        .Q(n359) );
  AO22X1 U382 ( .IN1(n2170), .IN2(wr_data[24]), .IN3(\r[9][24] ), .IN4(n2166),
        .Q(n360) );
  AO22X1 U383 ( .IN1(n2170), .IN2(wr_data[25]), .IN3(\r[9][25] ), .IN4(n2166),
        .Q(n361) );
  AO22X1 U384 ( .IN1(n2170), .IN2(wr_data[26]), .IN3(\r[9][26] ), .IN4(n2166),
        .Q(n362) );
  AO22X1 U385 ( .IN1(n2170), .IN2(wr_data[27]), .IN3(\r[9][27] ), .IN4(n2166),
        .Q(n363) );
  AO22X1 U386 ( .IN1(n2170), .IN2(wr_data[28]), .IN3(\r[9][28] ), .IN4(n2166),
        .Q(n364) );
  AO22X1 U387 ( .IN1(n2170), .IN2(wr_data[29]), .IN3(\r[9][29] ), .IN4(n2166),
        .Q(n365) );
  AO22X1 U388 ( .IN1(n2170), .IN2(wr_data[30]), .IN3(\r[9][30] ), .IN4(n2166),
        .Q(n366) );
  AO22X1 U389 ( .IN1(n2170), .IN2(wr_data[31]), .IN3(\r[9][31] ), .IN4(n2166),
        .Q(n367) );
  AO22X1 U390 ( .IN1(n2163), .IN2(wr_data[0]), .IN3(\r[10][0] ), .IN4(n56),
        .Q(n368) );
  AO22X1 U391 ( .IN1(n2163), .IN2(wr_data[1]), .IN3(\r[10][1] ), .IN4(n56),
        .Q(n369) );
  AO22X1 U392 ( .IN1(n2163), .IN2(wr_data[2]), .IN3(\r[10][2] ), .IN4(n56),
        .Q(n370) );
  AO22X1 U393 ( .IN1(n2163), .IN2(wr_data[3]), .IN3(\r[10][3] ), .IN4(n56),
        .Q(n371) );
  AO22X1 U394 ( .IN1(n2163), .IN2(wr_data[4]), .IN3(\r[10][4] ), .IN4(n56),
        .Q(n372) );
  AO22X1 U395 ( .IN1(n2163), .IN2(wr_data[5]), .IN3(\r[10][5] ), .IN4(n56),
        .Q(n373) );
  AO22X1 U396 ( .IN1(n2163), .IN2(wr_data[6]), .IN3(\r[10][6] ), .IN4(n56),
        .Q(n374) );
  AO22X1 U397 ( .IN1(n2163), .IN2(wr_data[7]), .IN3(\r[10][7] ), .IN4(n56),
        .Q(n375) );
  AO22X1 U398 ( .IN1(n2163), .IN2(wr_data[8]), .IN3(\r[10][8] ), .IN4(n2162),
        .Q(n376) );
  AO22X1 U399 ( .IN1(n2163), .IN2(wr_data[9]), .IN3(\r[10][9] ), .IN4(n2162),
        .Q(n377) );
  AO22X1 U400 ( .IN1(n2164), .IN2(wr_data[10]), .IN3(\r[10][10] ), .IN4(n2162),
        .Q(n378) );
  AO22X1 U401 ( .IN1(n2164), .IN2(wr_data[11]), .IN3(\r[10][11] ), .IN4(n2162),
        .Q(n379) );
  AO22X1 U402 ( .IN1(n2164), .IN2(wr_data[12]), .IN3(\r[10][12] ), .IN4(n2162),
        .Q(n380) );
  AO22X1 U403 ( .IN1(n2164), .IN2(wr_data[13]), .IN3(\r[10][13] ), .IN4(n2162),
        .Q(n381) );
  AO22X1 U404 ( .IN1(n2164), .IN2(wr_data[14]), .IN3(\r[10][14] ), .IN4(n2162),
        .Q(n382) );
  AO22X1 U405 ( .IN1(n2164), .IN2(wr_data[15]), .IN3(\r[10][15] ), .IN4(n2162),
        .Q(n383) );
  AO22X1 U406 ( .IN1(n2164), .IN2(wr_data[16]), .IN3(\r[10][16] ), .IN4(n2162),
        .Q(n384) );
  AO22X1 U407 ( .IN1(n2164), .IN2(wr_data[17]), .IN3(\r[10][17] ), .IN4(n2162),
        .Q(n385) );
  AO22X1 U408 ( .IN1(n2164), .IN2(wr_data[18]), .IN3(\r[10][18] ), .IN4(n2162),
        .Q(n386) );
  AO22X1 U409 ( .IN1(n2164), .IN2(wr_data[19]), .IN3(\r[10][19] ), .IN4(n2162),
        .Q(n387) );
  AO22X1 U410 ( .IN1(n2164), .IN2(wr_data[20]), .IN3(\r[10][20] ), .IN4(n2161),
        .Q(n388) );
  AO22X1 U411 ( .IN1(n2164), .IN2(wr_data[21]), .IN3(\r[10][21] ), .IN4(n2161),
        .Q(n389) );
  AO22X1 U412 ( .IN1(n2164), .IN2(wr_data[22]), .IN3(\r[10][22] ), .IN4(n2161),
        .Q(n390) );
  AO22X1 U413 ( .IN1(n2165), .IN2(wr_data[23]), .IN3(\r[10][23] ), .IN4(n2161),
        .Q(n391) );
  AO22X1 U414 ( .IN1(n2165), .IN2(wr_data[24]), .IN3(\r[10][24] ), .IN4(n2161),
        .Q(n392) );
  AO22X1 U415 ( .IN1(n2165), .IN2(wr_data[25]), .IN3(\r[10][25] ), .IN4(n2161),
        .Q(n393) );
  AO22X1 U416 ( .IN1(n2165), .IN2(wr_data[26]), .IN3(\r[10][26] ), .IN4(n2161),
        .Q(n394) );
  AO22X1 U417 ( .IN1(n2165), .IN2(wr_data[27]), .IN3(\r[10][27] ), .IN4(n2161),
        .Q(n395) );
  AO22X1 U418 ( .IN1(n2165), .IN2(wr_data[28]), .IN3(\r[10][28] ), .IN4(n2161),
        .Q(n396) );
  AO22X1 U419 ( .IN1(n2165), .IN2(wr_data[29]), .IN3(\r[10][29] ), .IN4(n2161),
        .Q(n397) );
  AO22X1 U420 ( .IN1(n2165), .IN2(wr_data[30]), .IN3(\r[10][30] ), .IN4(n2161),
        .Q(n398) );
  AO22X1 U421 ( .IN1(n2165), .IN2(wr_data[31]), .IN3(\r[10][31] ), .IN4(n2161),
        .Q(n399) );
  AO22X1 U422 ( .IN1(n2158), .IN2(wr_data[0]), .IN3(\r[11][0] ), .IN4(n57),
        .Q(n400) );
  AO22X1 U423 ( .IN1(n2158), .IN2(wr_data[1]), .IN3(\r[11][1] ), .IN4(n57),
        .Q(n401) );
  AO22X1 U424 ( .IN1(n2158), .IN2(wr_data[2]), .IN3(\r[11][2] ), .IN4(n57),
        .Q(n402) );
  AO22X1 U425 ( .IN1(n2158), .IN2(wr_data[3]), .IN3(\r[11][3] ), .IN4(n57),
        .Q(n403) );
  AO22X1 U426 ( .IN1(n2158), .IN2(wr_data[4]), .IN3(\r[11][4] ), .IN4(n57),
        .Q(n404) );
  AO22X1 U427 ( .IN1(n2158), .IN2(wr_data[5]), .IN3(\r[11][5] ), .IN4(n57),
        .Q(n405) );
  AO22X1 U428 ( .IN1(n2158), .IN2(wr_data[6]), .IN3(\r[11][6] ), .IN4(n57),
        .Q(n406) );
  AO22X1 U429 ( .IN1(n2158), .IN2(wr_data[7]), .IN3(\r[11][7] ), .IN4(n57),
        .Q(n407) );
  AO22X1 U430 ( .IN1(n2158), .IN2(wr_data[8]), .IN3(\r[11][8] ), .IN4(n2157),
        .Q(n408) );
  AO22X1 U431 ( .IN1(n2158), .IN2(wr_data[9]), .IN3(\r[11][9] ), .IN4(n2157),
        .Q(n409) );
  AO22X1 U432 ( .IN1(n2159), .IN2(wr_data[10]), .IN3(\r[11][10] ), .IN4(n2157),
        .Q(n410) );
  AO22X1 U433 ( .IN1(n2159), .IN2(wr_data[11]), .IN3(\r[11][11] ), .IN4(n2157),
        .Q(n411) );
  AO22X1 U434 ( .IN1(n2159), .IN2(wr_data[12]), .IN3(\r[11][12] ), .IN4(n2157),
        .Q(n412) );
  AO22X1 U435 ( .IN1(n2159), .IN2(wr_data[13]), .IN3(\r[11][13] ), .IN4(n2157),
        .Q(n413) );
  AO22X1 U436 ( .IN1(n2159), .IN2(wr_data[14]), .IN3(\r[11][14] ), .IN4(n2157),
        .Q(n414) );
  AO22X1 U437 ( .IN1(n2159), .IN2(wr_data[15]), .IN3(\r[11][15] ), .IN4(n2157),
        .Q(n415) );
  AO22X1 U438 ( .IN1(n2159), .IN2(wr_data[16]), .IN3(\r[11][16] ), .IN4(n2157),
        .Q(n416) );
  AO22X1 U439 ( .IN1(n2159), .IN2(wr_data[17]), .IN3(\r[11][17] ), .IN4(n2157),
        .Q(n417) );
  AO22X1 U440 ( .IN1(n2159), .IN2(wr_data[18]), .IN3(\r[11][18] ), .IN4(n2157),
        .Q(n418) );
  AO22X1 U441 ( .IN1(n2159), .IN2(wr_data[19]), .IN3(\r[11][19] ), .IN4(n2157),
        .Q(n419) );
  AO22X1 U442 ( .IN1(n2159), .IN2(wr_data[20]), .IN3(\r[11][20] ), .IN4(n2156),
        .Q(n420) );
  AO22X1 U443 ( .IN1(n2159), .IN2(wr_data[21]), .IN3(\r[11][21] ), .IN4(n2156),
        .Q(n421) );
  AO22X1 U444 ( .IN1(n2159), .IN2(wr_data[22]), .IN3(\r[11][22] ), .IN4(n2156),
        .Q(n422) );
  AO22X1 U445 ( .IN1(n2160), .IN2(wr_data[23]), .IN3(\r[11][23] ), .IN4(n2156),
        .Q(n423) );
  AO22X1 U446 ( .IN1(n2160), .IN2(wr_data[24]), .IN3(\r[11][24] ), .IN4(n2156),
        .Q(n424) );
  AO22X1 U447 ( .IN1(n2160), .IN2(wr_data[25]), .IN3(\r[11][25] ), .IN4(n2156),
        .Q(n425) );
  AO22X1 U448 ( .IN1(n2160), .IN2(wr_data[26]), .IN3(\r[11][26] ), .IN4(n2156),
        .Q(n426) );
  AO22X1 U449 ( .IN1(n2160), .IN2(wr_data[27]), .IN3(\r[11][27] ), .IN4(n2156),
        .Q(n427) );
  AO22X1 U450 ( .IN1(n2160), .IN2(wr_data[28]), .IN3(\r[11][28] ), .IN4(n2156),
        .Q(n428) );
  AO22X1 U451 ( .IN1(n2160), .IN2(wr_data[29]), .IN3(\r[11][29] ), .IN4(n2156),
        .Q(n429) );
  AO22X1 U452 ( .IN1(n2160), .IN2(wr_data[30]), .IN3(\r[11][30] ), .IN4(n2156),
        .Q(n430) );
  AO22X1 U453 ( .IN1(n2160), .IN2(wr_data[31]), .IN3(\r[11][31] ), .IN4(n2156),
        .Q(n431) );
  AO22X1 U454 ( .IN1(n2153), .IN2(wr_data[0]), .IN3(\r[12][0] ), .IN4(n58),
        .Q(n432) );
  AO22X1 U455 ( .IN1(n2153), .IN2(wr_data[1]), .IN3(\r[12][1] ), .IN4(n58),
        .Q(n433) );
  AO22X1 U456 ( .IN1(n2153), .IN2(wr_data[2]), .IN3(\r[12][2] ), .IN4(n58),
        .Q(n434) );
  AO22X1 U457 ( .IN1(n2153), .IN2(wr_data[3]), .IN3(\r[12][3] ), .IN4(n58),
        .Q(n435) );
  AO22X1 U458 ( .IN1(n2153), .IN2(wr_data[4]), .IN3(\r[12][4] ), .IN4(n58),
        .Q(n436) );
  AO22X1 U459 ( .IN1(n2153), .IN2(wr_data[5]), .IN3(\r[12][5] ), .IN4(n58),
        .Q(n437) );
  AO22X1 U460 ( .IN1(n2153), .IN2(wr_data[6]), .IN3(\r[12][6] ), .IN4(n58),
        .Q(n438) );
  AO22X1 U461 ( .IN1(n2153), .IN2(wr_data[7]), .IN3(\r[12][7] ), .IN4(n58),
        .Q(n439) );
  AO22X1 U462 ( .IN1(n2153), .IN2(wr_data[8]), .IN3(\r[12][8] ), .IN4(n2152),
        .Q(n440) );
  AO22X1 U463 ( .IN1(n2153), .IN2(wr_data[9]), .IN3(\r[12][9] ), .IN4(n2152),
        .Q(n441) );
  AO22X1 U464 ( .IN1(n2154), .IN2(wr_data[10]), .IN3(\r[12][10] ), .IN4(n2152),
        .Q(n442) );
  AO22X1 U465 ( .IN1(n2154), .IN2(wr_data[11]), .IN3(\r[12][11] ), .IN4(n2152),
        .Q(n443) );
  AO22X1 U466 ( .IN1(n2154), .IN2(wr_data[12]), .IN3(\r[12][12] ), .IN4(n2152),
        .Q(n444) );
  AO22X1 U467 ( .IN1(n2154), .IN2(wr_data[13]), .IN3(\r[12][13] ), .IN4(n2152),
        .Q(n445) );
  AO22X1 U468 ( .IN1(n2154), .IN2(wr_data[14]), .IN3(\r[12][14] ), .IN4(n2152),
        .Q(n446) );
  AO22X1 U469 ( .IN1(n2154), .IN2(wr_data[15]), .IN3(\r[12][15] ), .IN4(n2152),
        .Q(n447) );
  AO22X1 U470 ( .IN1(n2154), .IN2(wr_data[16]), .IN3(\r[12][16] ), .IN4(n2152),
        .Q(n448) );
  AO22X1 U471 ( .IN1(n2154), .IN2(wr_data[17]), .IN3(\r[12][17] ), .IN4(n2152),
        .Q(n449) );
  AO22X1 U472 ( .IN1(n2154), .IN2(wr_data[18]), .IN3(\r[12][18] ), .IN4(n2152),
        .Q(n450) );
  AO22X1 U473 ( .IN1(n2154), .IN2(wr_data[19]), .IN3(\r[12][19] ), .IN4(n2152),
        .Q(n451) );
  AO22X1 U474 ( .IN1(n2154), .IN2(wr_data[20]), .IN3(\r[12][20] ), .IN4(n2151),
        .Q(n452) );
  AO22X1 U475 ( .IN1(n2154), .IN2(wr_data[21]), .IN3(\r[12][21] ), .IN4(n2151),
        .Q(n453) );
  AO22X1 U476 ( .IN1(n2154), .IN2(wr_data[22]), .IN3(\r[12][22] ), .IN4(n2151),
        .Q(n454) );
  AO22X1 U477 ( .IN1(n2155), .IN2(wr_data[23]), .IN3(\r[12][23] ), .IN4(n2151),
        .Q(n455) );
  AO22X1 U478 ( .IN1(n2155), .IN2(wr_data[24]), .IN3(\r[12][24] ), .IN4(n2151),
        .Q(n456) );
  AO22X1 U479 ( .IN1(n2155), .IN2(wr_data[25]), .IN3(\r[12][25] ), .IN4(n2151),
        .Q(n457) );
  AO22X1 U480 ( .IN1(n2155), .IN2(wr_data[26]), .IN3(\r[12][26] ), .IN4(n2151),
        .Q(n458) );
  AO22X1 U481 ( .IN1(n2155), .IN2(wr_data[27]), .IN3(\r[12][27] ), .IN4(n2151),
        .Q(n459) );
  AO22X1 U482 ( .IN1(n2155), .IN2(wr_data[28]), .IN3(\r[12][28] ), .IN4(n2151),
        .Q(n460) );
  AO22X1 U483 ( .IN1(n2155), .IN2(wr_data[29]), .IN3(\r[12][29] ), .IN4(n2151),
        .Q(n461) );
  AO22X1 U484 ( .IN1(n2155), .IN2(wr_data[30]), .IN3(\r[12][30] ), .IN4(n2151),
        .Q(n462) );
  AO22X1 U485 ( .IN1(n2155), .IN2(wr_data[31]), .IN3(\r[12][31] ), .IN4(n2151),
        .Q(n463) );
  AO22X1 U486 ( .IN1(n2148), .IN2(wr_data[0]), .IN3(\r[13][0] ), .IN4(n59),
        .Q(n464) );
  AO22X1 U487 ( .IN1(n2148), .IN2(wr_data[1]), .IN3(\r[13][1] ), .IN4(n59),
        .Q(n465) );
  AO22X1 U488 ( .IN1(n2148), .IN2(wr_data[2]), .IN3(\r[13][2] ), .IN4(n59),
        .Q(n466) );
  AO22X1 U489 ( .IN1(n2148), .IN2(wr_data[3]), .IN3(\r[13][3] ), .IN4(n59),
        .Q(n467) );
  AO22X1 U490 ( .IN1(n2148), .IN2(wr_data[4]), .IN3(\r[13][4] ), .IN4(n59),
        .Q(n468) );
  AO22X1 U491 ( .IN1(n2148), .IN2(wr_data[5]), .IN3(\r[13][5] ), .IN4(n59),
        .Q(n469) );
  AO22X1 U492 ( .IN1(n2148), .IN2(wr_data[6]), .IN3(\r[13][6] ), .IN4(n59),
        .Q(n470) );
  AO22X1 U493 ( .IN1(n2148), .IN2(wr_data[7]), .IN3(\r[13][7] ), .IN4(n59),
        .Q(n471) );
  AO22X1 U494 ( .IN1(n2148), .IN2(wr_data[8]), .IN3(\r[13][8] ), .IN4(n2147),
        .Q(n472) );
  AO22X1 U495 ( .IN1(n2148), .IN2(wr_data[9]), .IN3(\r[13][9] ), .IN4(n2147),
        .Q(n473) );
  AO22X1 U496 ( .IN1(n2149), .IN2(wr_data[10]), .IN3(\r[13][10] ), .IN4(n2147),
        .Q(n474) );
  AO22X1 U497 ( .IN1(n2149), .IN2(wr_data[11]), .IN3(\r[13][11] ), .IN4(n2147),
        .Q(n475) );
  AO22X1 U498 ( .IN1(n2149), .IN2(wr_data[12]), .IN3(\r[13][12] ), .IN4(n2147),
        .Q(n476) );
  AO22X1 U499 ( .IN1(n2149), .IN2(wr_data[13]), .IN3(\r[13][13] ), .IN4(n2147),
        .Q(n477) );
  AO22X1 U500 ( .IN1(n2149), .IN2(wr_data[14]), .IN3(\r[13][14] ), .IN4(n2147),
        .Q(n478) );
  AO22X1 U501 ( .IN1(n2149), .IN2(wr_data[15]), .IN3(\r[13][15] ), .IN4(n2147),
        .Q(n479) );
  AO22X1 U502 ( .IN1(n2149), .IN2(wr_data[16]), .IN3(\r[13][16] ), .IN4(n2147),
        .Q(n480) );
  AO22X1 U503 ( .IN1(n2149), .IN2(wr_data[17]), .IN3(\r[13][17] ), .IN4(n2147),
        .Q(n481) );
  AO22X1 U504 ( .IN1(n2149), .IN2(wr_data[18]), .IN3(\r[13][18] ), .IN4(n2147),
        .Q(n482) );
  AO22X1 U505 ( .IN1(n2149), .IN2(wr_data[19]), .IN3(\r[13][19] ), .IN4(n2147),
        .Q(n483) );
  AO22X1 U506 ( .IN1(n2149), .IN2(wr_data[20]), .IN3(\r[13][20] ), .IN4(n2146),
        .Q(n484) );
  AO22X1 U507 ( .IN1(n2149), .IN2(wr_data[21]), .IN3(\r[13][21] ), .IN4(n2146),
        .Q(n485) );
  AO22X1 U508 ( .IN1(n2149), .IN2(wr_data[22]), .IN3(\r[13][22] ), .IN4(n2146),
        .Q(n486) );
  AO22X1 U509 ( .IN1(n2150), .IN2(wr_data[23]), .IN3(\r[13][23] ), .IN4(n2146),
        .Q(n487) );
  AO22X1 U510 ( .IN1(n2150), .IN2(wr_data[24]), .IN3(\r[13][24] ), .IN4(n2146),
        .Q(n488) );
  AO22X1 U511 ( .IN1(n2150), .IN2(wr_data[25]), .IN3(\r[13][25] ), .IN4(n2146),
        .Q(n489) );
  AO22X1 U512 ( .IN1(n2150), .IN2(wr_data[26]), .IN3(\r[13][26] ), .IN4(n2146),
        .Q(n490) );
  AO22X1 U513 ( .IN1(n2150), .IN2(wr_data[27]), .IN3(\r[13][27] ), .IN4(n2146),
        .Q(n491) );
  AO22X1 U514 ( .IN1(n2150), .IN2(wr_data[28]), .IN3(\r[13][28] ), .IN4(n2146),
        .Q(n492) );
  AO22X1 U515 ( .IN1(n2150), .IN2(wr_data[29]), .IN3(\r[13][29] ), .IN4(n2146),
        .Q(n493) );
  AO22X1 U516 ( .IN1(n2150), .IN2(wr_data[30]), .IN3(\r[13][30] ), .IN4(n2146),
        .Q(n494) );
  AO22X1 U517 ( .IN1(n2150), .IN2(wr_data[31]), .IN3(\r[13][31] ), .IN4(n2146),
        .Q(n495) );
  AO22X1 U518 ( .IN1(n2143), .IN2(wr_data[0]), .IN3(\r[14][0] ), .IN4(n60),
        .Q(n496) );
  AO22X1 U519 ( .IN1(n2143), .IN2(wr_data[1]), .IN3(\r[14][1] ), .IN4(n60),
        .Q(n497) );
  AO22X1 U520 ( .IN1(n2143), .IN2(wr_data[2]), .IN3(\r[14][2] ), .IN4(n60),
        .Q(n498) );
  AO22X1 U521 ( .IN1(n2143), .IN2(wr_data[3]), .IN3(\r[14][3] ), .IN4(n60),
        .Q(n499) );
  AO22X1 U522 ( .IN1(n2143), .IN2(wr_data[4]), .IN3(\r[14][4] ), .IN4(n60),
        .Q(n500) );
  AO22X1 U523 ( .IN1(n2143), .IN2(wr_data[5]), .IN3(\r[14][5] ), .IN4(n60),
        .Q(n501) );
  AO22X1 U524 ( .IN1(n2143), .IN2(wr_data[6]), .IN3(\r[14][6] ), .IN4(n60),
        .Q(n502) );
  AO22X1 U525 ( .IN1(n2143), .IN2(wr_data[7]), .IN3(\r[14][7] ), .IN4(n60),
        .Q(n503) );
  AO22X1 U526 ( .IN1(n2143), .IN2(wr_data[8]), .IN3(\r[14][8] ), .IN4(n2142),
        .Q(n504) );
  AO22X1 U527 ( .IN1(n2143), .IN2(wr_data[9]), .IN3(\r[14][9] ), .IN4(n2142),
        .Q(n505) );
  AO22X1 U528 ( .IN1(n2144), .IN2(wr_data[10]), .IN3(\r[14][10] ), .IN4(n2142),
        .Q(n506) );
  AO22X1 U529 ( .IN1(n2144), .IN2(wr_data[11]), .IN3(\r[14][11] ), .IN4(n2142),
        .Q(n507) );
  AO22X1 U530 ( .IN1(n2144), .IN2(wr_data[12]), .IN3(\r[14][12] ), .IN4(n2142),
        .Q(n508) );
  AO22X1 U531 ( .IN1(n2144), .IN2(wr_data[13]), .IN3(\r[14][13] ), .IN4(n2142),
        .Q(n509) );
  AO22X1 U532 ( .IN1(n2144), .IN2(wr_data[14]), .IN3(\r[14][14] ), .IN4(n2142),
        .Q(n510) );
  AO22X1 U533 ( .IN1(n2144), .IN2(wr_data[15]), .IN3(\r[14][15] ), .IN4(n2142),
        .Q(n511) );
  AO22X1 U534 ( .IN1(n2144), .IN2(wr_data[16]), .IN3(\r[14][16] ), .IN4(n2142),
        .Q(n512) );
  AO22X1 U535 ( .IN1(n2144), .IN2(wr_data[17]), .IN3(\r[14][17] ), .IN4(n2142),
        .Q(n513) );
  AO22X1 U536 ( .IN1(n2144), .IN2(wr_data[18]), .IN3(\r[14][18] ), .IN4(n2142),
        .Q(n514) );
  AO22X1 U537 ( .IN1(n2144), .IN2(wr_data[19]), .IN3(\r[14][19] ), .IN4(n2142),
        .Q(n515) );
  AO22X1 U538 ( .IN1(n2144), .IN2(wr_data[20]), .IN3(\r[14][20] ), .IN4(n2141),
        .Q(n516) );
  AO22X1 U539 ( .IN1(n2144), .IN2(wr_data[21]), .IN3(\r[14][21] ), .IN4(n2141),
        .Q(n517) );
  AO22X1 U540 ( .IN1(n2144), .IN2(wr_data[22]), .IN3(\r[14][22] ), .IN4(n2141),
        .Q(n518) );
  AO22X1 U541 ( .IN1(n2145), .IN2(wr_data[23]), .IN3(\r[14][23] ), .IN4(n2141),
        .Q(n519) );
  AO22X1 U542 ( .IN1(n2145), .IN2(wr_data[24]), .IN3(\r[14][24] ), .IN4(n2141),
        .Q(n520) );
  AO22X1 U543 ( .IN1(n2145), .IN2(wr_data[25]), .IN3(\r[14][25] ), .IN4(n2141),
        .Q(n521) );
  AO22X1 U544 ( .IN1(n2145), .IN2(wr_data[26]), .IN3(\r[14][26] ), .IN4(n2141),
        .Q(n522) );
  AO22X1 U545 ( .IN1(n2145), .IN2(wr_data[27]), .IN3(\r[14][27] ), .IN4(n2141),
        .Q(n523) );
  AO22X1 U546 ( .IN1(n2145), .IN2(wr_data[28]), .IN3(\r[14][28] ), .IN4(n2141),
        .Q(n524) );
  AO22X1 U547 ( .IN1(n2145), .IN2(wr_data[29]), .IN3(\r[14][29] ), .IN4(n2141),
        .Q(n525) );
  AO22X1 U548 ( .IN1(n2145), .IN2(wr_data[30]), .IN3(\r[14][30] ), .IN4(n2141),
        .Q(n526) );
  AO22X1 U549 ( .IN1(n2145), .IN2(wr_data[31]), .IN3(\r[14][31] ), .IN4(n2141),
        .Q(n527) );
  AO22X1 U550 ( .IN1(n2138), .IN2(wr_data[0]), .IN3(\r[15][0] ), .IN4(n61),
        .Q(n528) );
  AO22X1 U551 ( .IN1(n2138), .IN2(wr_data[1]), .IN3(\r[15][1] ), .IN4(n61),
        .Q(n529) );
  AO22X1 U552 ( .IN1(n2138), .IN2(wr_data[2]), .IN3(\r[15][2] ), .IN4(n61),
        .Q(n530) );
  AO22X1 U553 ( .IN1(n2138), .IN2(wr_data[3]), .IN3(\r[15][3] ), .IN4(n61),
        .Q(n531) );
  AO22X1 U554 ( .IN1(n2138), .IN2(wr_data[4]), .IN3(\r[15][4] ), .IN4(n61),
        .Q(n532) );
  AO22X1 U555 ( .IN1(n2138), .IN2(wr_data[5]), .IN3(\r[15][5] ), .IN4(n61),
        .Q(n533) );
  AO22X1 U556 ( .IN1(n2138), .IN2(wr_data[6]), .IN3(\r[15][6] ), .IN4(n61),
        .Q(n534) );
  AO22X1 U557 ( .IN1(n2138), .IN2(wr_data[7]), .IN3(\r[15][7] ), .IN4(n61),
        .Q(n535) );
  AO22X1 U558 ( .IN1(n2138), .IN2(wr_data[8]), .IN3(\r[15][8] ), .IN4(n2137),
        .Q(n536) );
  AO22X1 U559 ( .IN1(n2138), .IN2(wr_data[9]), .IN3(\r[15][9] ), .IN4(n2137),
        .Q(n537) );
  AO22X1 U560 ( .IN1(n2139), .IN2(wr_data[10]), .IN3(\r[15][10] ), .IN4(n2137),
        .Q(n538) );
  AO22X1 U561 ( .IN1(n2139), .IN2(wr_data[11]), .IN3(\r[15][11] ), .IN4(n2137),
        .Q(n539) );
  AO22X1 U562 ( .IN1(n2139), .IN2(wr_data[12]), .IN3(\r[15][12] ), .IN4(n2137),
        .Q(n540) );
  AO22X1 U563 ( .IN1(n2139), .IN2(wr_data[13]), .IN3(\r[15][13] ), .IN4(n2137),
        .Q(n541) );
  AO22X1 U564 ( .IN1(n2139), .IN2(wr_data[14]), .IN3(\r[15][14] ), .IN4(n2137),
        .Q(n542) );
  AO22X1 U565 ( .IN1(n2139), .IN2(wr_data[15]), .IN3(\r[15][15] ), .IN4(n2137),
        .Q(n543) );
  AO22X1 U566 ( .IN1(n2139), .IN2(wr_data[16]), .IN3(\r[15][16] ), .IN4(n2137),
        .Q(n544) );
  AO22X1 U567 ( .IN1(n2139), .IN2(wr_data[17]), .IN3(\r[15][17] ), .IN4(n2137),
        .Q(n545) );
  AO22X1 U568 ( .IN1(n2139), .IN2(wr_data[18]), .IN3(\r[15][18] ), .IN4(n2137),
        .Q(n546) );
  AO22X1 U569 ( .IN1(n2139), .IN2(wr_data[19]), .IN3(\r[15][19] ), .IN4(n2137),
        .Q(n547) );
  AO22X1 U570 ( .IN1(n2139), .IN2(wr_data[20]), .IN3(\r[15][20] ), .IN4(n2136),
        .Q(n548) );
  AO22X1 U571 ( .IN1(n2139), .IN2(wr_data[21]), .IN3(\r[15][21] ), .IN4(n2136),
        .Q(n549) );
  AO22X1 U572 ( .IN1(n2139), .IN2(wr_data[22]), .IN3(\r[15][22] ), .IN4(n2136),
        .Q(n550) );
  AO22X1 U573 ( .IN1(n2140), .IN2(wr_data[23]), .IN3(\r[15][23] ), .IN4(n2136),
        .Q(n551) );
  AO22X1 U574 ( .IN1(n2140), .IN2(wr_data[24]), .IN3(\r[15][24] ), .IN4(n2136),
        .Q(n552) );
  AO22X1 U575 ( .IN1(n2140), .IN2(wr_data[25]), .IN3(\r[15][25] ), .IN4(n2136),
        .Q(n553) );
  AO22X1 U576 ( .IN1(n2140), .IN2(wr_data[26]), .IN3(\r[15][26] ), .IN4(n2136),
        .Q(n554) );
  AO22X1 U577 ( .IN1(n2140), .IN2(wr_data[27]), .IN3(\r[15][27] ), .IN4(n2136),
        .Q(n555) );
  AO22X1 U578 ( .IN1(n2140), .IN2(wr_data[28]), .IN3(\r[15][28] ), .IN4(n2136),
        .Q(n556) );
  AO22X1 U579 ( .IN1(n2140), .IN2(wr_data[29]), .IN3(\r[15][29] ), .IN4(n2136),
        .Q(n557) );
  AO22X1 U580 ( .IN1(n2140), .IN2(wr_data[30]), .IN3(\r[15][30] ), .IN4(n2136),
        .Q(n558) );
  AO22X1 U581 ( .IN1(n2140), .IN2(wr_data[31]), .IN3(\r[15][31] ), .IN4(n2136),
        .Q(n559) );
  AND3X1 U582 ( .IN1(wr_en), .IN2(n2299), .IN3(wr_addr[3]), .Q(n54) );
  AO22X1 U583 ( .IN1(n2133), .IN2(wr_data[0]), .IN3(\r[16][0] ), .IN4(n62),
        .Q(n560) );
  AO22X1 U584 ( .IN1(n2133), .IN2(wr_data[1]), .IN3(\r[16][1] ), .IN4(n62),
        .Q(n561) );
  AO22X1 U585 ( .IN1(n2133), .IN2(wr_data[2]), .IN3(\r[16][2] ), .IN4(n62),
        .Q(n562) );
  AO22X1 U586 ( .IN1(n2133), .IN2(wr_data[3]), .IN3(\r[16][3] ), .IN4(n62),
        .Q(n563) );
  AO22X1 U587 ( .IN1(n2133), .IN2(wr_data[4]), .IN3(\r[16][4] ), .IN4(n62),
        .Q(n564) );
  AO22X1 U588 ( .IN1(n2133), .IN2(wr_data[5]), .IN3(\r[16][5] ), .IN4(n62),
        .Q(n565) );
  AO22X1 U589 ( .IN1(n2133), .IN2(wr_data[6]), .IN3(\r[16][6] ), .IN4(n62),
        .Q(n566) );
  AO22X1 U590 ( .IN1(n2133), .IN2(wr_data[7]), .IN3(\r[16][7] ), .IN4(n62),
        .Q(n567) );
  AO22X1 U591 ( .IN1(n2133), .IN2(wr_data[8]), .IN3(\r[16][8] ), .IN4(n2132),
        .Q(n568) );
  AO22X1 U592 ( .IN1(n2133), .IN2(wr_data[9]), .IN3(\r[16][9] ), .IN4(n2132),
        .Q(n569) );
  AO22X1 U593 ( .IN1(n2134), .IN2(wr_data[10]), .IN3(\r[16][10] ), .IN4(n2132),
        .Q(n570) );
  AO22X1 U594 ( .IN1(n2134), .IN2(wr_data[11]), .IN3(\r[16][11] ), .IN4(n2132),
        .Q(n571) );
  AO22X1 U595 ( .IN1(n2134), .IN2(wr_data[12]), .IN3(\r[16][12] ), .IN4(n2132),
        .Q(n572) );
  AO22X1 U596 ( .IN1(n2134), .IN2(wr_data[13]), .IN3(\r[16][13] ), .IN4(n2132),
        .Q(n573) );
  AO22X1 U597 ( .IN1(n2134), .IN2(wr_data[14]), .IN3(\r[16][14] ), .IN4(n2132),
        .Q(n574) );
  AO22X1 U598 ( .IN1(n2134), .IN2(wr_data[15]), .IN3(\r[16][15] ), .IN4(n2132),
        .Q(n575) );
  AO22X1 U599 ( .IN1(n2134), .IN2(wr_data[16]), .IN3(\r[16][16] ), .IN4(n2132),
        .Q(n576) );
  AO22X1 U600 ( .IN1(n2134), .IN2(wr_data[17]), .IN3(\r[16][17] ), .IN4(n2132),
        .Q(n577) );
  AO22X1 U601 ( .IN1(n2134), .IN2(wr_data[18]), .IN3(\r[16][18] ), .IN4(n2132),
        .Q(n578) );
  AO22X1 U602 ( .IN1(n2134), .IN2(wr_data[19]), .IN3(\r[16][19] ), .IN4(n2132),
        .Q(n579) );
  AO22X1 U603 ( .IN1(n2134), .IN2(wr_data[20]), .IN3(\r[16][20] ), .IN4(n2131),
        .Q(n580) );
  AO22X1 U604 ( .IN1(n2134), .IN2(wr_data[21]), .IN3(\r[16][21] ), .IN4(n2131),
        .Q(n581) );
  AO22X1 U605 ( .IN1(n2134), .IN2(wr_data[22]), .IN3(\r[16][22] ), .IN4(n2131),
        .Q(n582) );
  AO22X1 U606 ( .IN1(n2135), .IN2(wr_data[23]), .IN3(\r[16][23] ), .IN4(n2131),
        .Q(n583) );
  AO22X1 U607 ( .IN1(n2135), .IN2(wr_data[24]), .IN3(\r[16][24] ), .IN4(n2131),
        .Q(n584) );
  AO22X1 U608 ( .IN1(n2135), .IN2(wr_data[25]), .IN3(\r[16][25] ), .IN4(n2131),
        .Q(n585) );
  AO22X1 U609 ( .IN1(n2135), .IN2(wr_data[26]), .IN3(\r[16][26] ), .IN4(n2131),
        .Q(n586) );
  AO22X1 U610 ( .IN1(n2135), .IN2(wr_data[27]), .IN3(\r[16][27] ), .IN4(n2131),
        .Q(n587) );
  AO22X1 U611 ( .IN1(n2135), .IN2(wr_data[28]), .IN3(\r[16][28] ), .IN4(n2131),
        .Q(n588) );
  AO22X1 U612 ( .IN1(n2135), .IN2(wr_data[29]), .IN3(\r[16][29] ), .IN4(n2131),
        .Q(n589) );
  AO22X1 U613 ( .IN1(n2135), .IN2(wr_data[30]), .IN3(\r[16][30] ), .IN4(n2131),
        .Q(n590) );
  AO22X1 U614 ( .IN1(n2135), .IN2(wr_data[31]), .IN3(\r[16][31] ), .IN4(n2131),
        .Q(n591) );
  AO22X1 U615 ( .IN1(n2128), .IN2(wr_data[0]), .IN3(\r[17][0] ), .IN4(n64),
        .Q(n592) );
  AO22X1 U616 ( .IN1(n2128), .IN2(wr_data[1]), .IN3(\r[17][1] ), .IN4(n64),
        .Q(n593) );
  AO22X1 U617 ( .IN1(n2128), .IN2(wr_data[2]), .IN3(\r[17][2] ), .IN4(n64),
        .Q(n594) );
  AO22X1 U618 ( .IN1(n2128), .IN2(wr_data[3]), .IN3(\r[17][3] ), .IN4(n64),
        .Q(n595) );
  AO22X1 U619 ( .IN1(n2128), .IN2(wr_data[4]), .IN3(\r[17][4] ), .IN4(n64),
        .Q(n596) );
  AO22X1 U620 ( .IN1(n2128), .IN2(wr_data[5]), .IN3(\r[17][5] ), .IN4(n64),
        .Q(n597) );
  AO22X1 U621 ( .IN1(n2128), .IN2(wr_data[6]), .IN3(\r[17][6] ), .IN4(n64),
        .Q(n598) );
  AO22X1 U622 ( .IN1(n2128), .IN2(wr_data[7]), .IN3(\r[17][7] ), .IN4(n64),
        .Q(n599) );
  AO22X1 U623 ( .IN1(n2128), .IN2(wr_data[8]), .IN3(\r[17][8] ), .IN4(n2127),
        .Q(n600) );
  AO22X1 U624 ( .IN1(n2128), .IN2(wr_data[9]), .IN3(\r[17][9] ), .IN4(n2127),
        .Q(n601) );
  AO22X1 U625 ( .IN1(n2129), .IN2(wr_data[10]), .IN3(\r[17][10] ), .IN4(n2127),
        .Q(n602) );
  AO22X1 U626 ( .IN1(n2129), .IN2(wr_data[11]), .IN3(\r[17][11] ), .IN4(n2127),
        .Q(n603) );
  AO22X1 U627 ( .IN1(n2129), .IN2(wr_data[12]), .IN3(\r[17][12] ), .IN4(n2127),
        .Q(n604) );
  AO22X1 U628 ( .IN1(n2129), .IN2(wr_data[13]), .IN3(\r[17][13] ), .IN4(n2127),
        .Q(n605) );
  AO22X1 U629 ( .IN1(n2129), .IN2(wr_data[14]), .IN3(\r[17][14] ), .IN4(n2127),
        .Q(n606) );
  AO22X1 U630 ( .IN1(n2129), .IN2(wr_data[15]), .IN3(\r[17][15] ), .IN4(n2127),
        .Q(n607) );
  AO22X1 U631 ( .IN1(n2129), .IN2(wr_data[16]), .IN3(\r[17][16] ), .IN4(n2127),
        .Q(n608) );
  AO22X1 U632 ( .IN1(n2129), .IN2(wr_data[17]), .IN3(\r[17][17] ), .IN4(n2127),
        .Q(n609) );
  AO22X1 U633 ( .IN1(n2129), .IN2(wr_data[18]), .IN3(\r[17][18] ), .IN4(n2127),
        .Q(n610) );
  AO22X1 U634 ( .IN1(n2129), .IN2(wr_data[19]), .IN3(\r[17][19] ), .IN4(n2127),
        .Q(n611) );
  AO22X1 U635 ( .IN1(n2129), .IN2(wr_data[20]), .IN3(\r[17][20] ), .IN4(n2126),
        .Q(n612) );
  AO22X1 U636 ( .IN1(n2129), .IN2(wr_data[21]), .IN3(\r[17][21] ), .IN4(n2126),
        .Q(n613) );
  AO22X1 U637 ( .IN1(n2129), .IN2(wr_data[22]), .IN3(\r[17][22] ), .IN4(n2126),
        .Q(n614) );
  AO22X1 U638 ( .IN1(n2130), .IN2(wr_data[23]), .IN3(\r[17][23] ), .IN4(n2126),
        .Q(n615) );
  AO22X1 U639 ( .IN1(n2130), .IN2(wr_data[24]), .IN3(\r[17][24] ), .IN4(n2126),
        .Q(n616) );
  AO22X1 U640 ( .IN1(n2130), .IN2(wr_data[25]), .IN3(\r[17][25] ), .IN4(n2126),
        .Q(n617) );
  AO22X1 U641 ( .IN1(n2130), .IN2(wr_data[26]), .IN3(\r[17][26] ), .IN4(n2126),
        .Q(n618) );
  AO22X1 U642 ( .IN1(n2130), .IN2(wr_data[27]), .IN3(\r[17][27] ), .IN4(n2126),
        .Q(n619) );
  AO22X1 U643 ( .IN1(n2130), .IN2(wr_data[28]), .IN3(\r[17][28] ), .IN4(n2126),
        .Q(n620) );
  AO22X1 U644 ( .IN1(n2130), .IN2(wr_data[29]), .IN3(\r[17][29] ), .IN4(n2126),
        .Q(n621) );
  AO22X1 U645 ( .IN1(n2130), .IN2(wr_data[30]), .IN3(\r[17][30] ), .IN4(n2126),
        .Q(n622) );
  AO22X1 U646 ( .IN1(n2130), .IN2(wr_data[31]), .IN3(\r[17][31] ), .IN4(n2126),
        .Q(n623) );
  AO22X1 U647 ( .IN1(n2123), .IN2(wr_data[0]), .IN3(\r[18][0] ), .IN4(n65),
        .Q(n624) );
  AO22X1 U648 ( .IN1(n2123), .IN2(wr_data[1]), .IN3(\r[18][1] ), .IN4(n65),
        .Q(n625) );
  AO22X1 U649 ( .IN1(n2123), .IN2(wr_data[2]), .IN3(\r[18][2] ), .IN4(n65),
        .Q(n626) );
  AO22X1 U650 ( .IN1(n2123), .IN2(wr_data[3]), .IN3(\r[18][3] ), .IN4(n65),
        .Q(n627) );
  AO22X1 U651 ( .IN1(n2123), .IN2(wr_data[4]), .IN3(\r[18][4] ), .IN4(n65),
        .Q(n628) );
  AO22X1 U652 ( .IN1(n2123), .IN2(wr_data[5]), .IN3(\r[18][5] ), .IN4(n65),
        .Q(n629) );
  AO22X1 U653 ( .IN1(n2123), .IN2(wr_data[6]), .IN3(\r[18][6] ), .IN4(n65),
        .Q(n630) );
  AO22X1 U654 ( .IN1(n2123), .IN2(wr_data[7]), .IN3(\r[18][7] ), .IN4(n65),
        .Q(n631) );
  AO22X1 U655 ( .IN1(n2123), .IN2(wr_data[8]), .IN3(\r[18][8] ), .IN4(n2122),
        .Q(n632) );
  AO22X1 U656 ( .IN1(n2123), .IN2(wr_data[9]), .IN3(\r[18][9] ), .IN4(n2122),
        .Q(n633) );
  AO22X1 U657 ( .IN1(n2124), .IN2(wr_data[10]), .IN3(\r[18][10] ), .IN4(n2122),
        .Q(n634) );
  AO22X1 U658 ( .IN1(n2124), .IN2(wr_data[11]), .IN3(\r[18][11] ), .IN4(n2122),
        .Q(n635) );
  AO22X1 U659 ( .IN1(n2124), .IN2(wr_data[12]), .IN3(\r[18][12] ), .IN4(n2122),
        .Q(n636) );
  AO22X1 U660 ( .IN1(n2124), .IN2(wr_data[13]), .IN3(\r[18][13] ), .IN4(n2122),
        .Q(n637) );
  AO22X1 U661 ( .IN1(n2124), .IN2(wr_data[14]), .IN3(\r[18][14] ), .IN4(n2122),
        .Q(n638) );
  AO22X1 U662 ( .IN1(n2124), .IN2(wr_data[15]), .IN3(\r[18][15] ), .IN4(n2122),
        .Q(n639) );
  AO22X1 U663 ( .IN1(n2124), .IN2(wr_data[16]), .IN3(\r[18][16] ), .IN4(n2122),
        .Q(n640) );
  AO22X1 U664 ( .IN1(n2124), .IN2(wr_data[17]), .IN3(\r[18][17] ), .IN4(n2122),
        .Q(n641) );
  AO22X1 U665 ( .IN1(n2124), .IN2(wr_data[18]), .IN3(\r[18][18] ), .IN4(n2122),
        .Q(n642) );
  AO22X1 U666 ( .IN1(n2124), .IN2(wr_data[19]), .IN3(\r[18][19] ), .IN4(n2122),
        .Q(n643) );
  AO22X1 U667 ( .IN1(n2124), .IN2(wr_data[20]), .IN3(\r[18][20] ), .IN4(n2121),
        .Q(n644) );
  AO22X1 U668 ( .IN1(n2124), .IN2(wr_data[21]), .IN3(\r[18][21] ), .IN4(n2121),
        .Q(n645) );
  AO22X1 U669 ( .IN1(n2124), .IN2(wr_data[22]), .IN3(\r[18][22] ), .IN4(n2121),
        .Q(n646) );
  AO22X1 U670 ( .IN1(n2125), .IN2(wr_data[23]), .IN3(\r[18][23] ), .IN4(n2121),
        .Q(n647) );
  AO22X1 U671 ( .IN1(n2125), .IN2(wr_data[24]), .IN3(\r[18][24] ), .IN4(n2121),
        .Q(n648) );
  AO22X1 U672 ( .IN1(n2125), .IN2(wr_data[25]), .IN3(\r[18][25] ), .IN4(n2121),
        .Q(n649) );
  AO22X1 U673 ( .IN1(n2125), .IN2(wr_data[26]), .IN3(\r[18][26] ), .IN4(n2121),
        .Q(n650) );
  AO22X1 U674 ( .IN1(n2125), .IN2(wr_data[27]), .IN3(\r[18][27] ), .IN4(n2121),
        .Q(n651) );
  AO22X1 U675 ( .IN1(n2125), .IN2(wr_data[28]), .IN3(\r[18][28] ), .IN4(n2121),
        .Q(n652) );
  AO22X1 U676 ( .IN1(n2125), .IN2(wr_data[29]), .IN3(\r[18][29] ), .IN4(n2121),
        .Q(n653) );
  AO22X1 U677 ( .IN1(n2125), .IN2(wr_data[30]), .IN3(\r[18][30] ), .IN4(n2121),
        .Q(n654) );
  AO22X1 U678 ( .IN1(n2125), .IN2(wr_data[31]), .IN3(\r[18][31] ), .IN4(n2121),
        .Q(n655) );
  AO22X1 U679 ( .IN1(n2118), .IN2(wr_data[0]), .IN3(\r[19][0] ), .IN4(n66),
        .Q(n656) );
  AO22X1 U680 ( .IN1(n2118), .IN2(wr_data[1]), .IN3(\r[19][1] ), .IN4(n66),
        .Q(n657) );
  AO22X1 U681 ( .IN1(n2118), .IN2(wr_data[2]), .IN3(\r[19][2] ), .IN4(n66),
        .Q(n658) );
  AO22X1 U682 ( .IN1(n2118), .IN2(wr_data[3]), .IN3(\r[19][3] ), .IN4(n66),
        .Q(n659) );
  AO22X1 U683 ( .IN1(n2118), .IN2(wr_data[4]), .IN3(\r[19][4] ), .IN4(n66),
        .Q(n660) );
  AO22X1 U684 ( .IN1(n2118), .IN2(wr_data[5]), .IN3(\r[19][5] ), .IN4(n66),
        .Q(n661) );
  AO22X1 U685 ( .IN1(n2118), .IN2(wr_data[6]), .IN3(\r[19][6] ), .IN4(n66),
        .Q(n662) );
  AO22X1 U686 ( .IN1(n2118), .IN2(wr_data[7]), .IN3(\r[19][7] ), .IN4(n66),
        .Q(n663) );
  AO22X1 U687 ( .IN1(n2118), .IN2(wr_data[8]), .IN3(\r[19][8] ), .IN4(n2117),
        .Q(n664) );
  AO22X1 U688 ( .IN1(n2118), .IN2(wr_data[9]), .IN3(\r[19][9] ), .IN4(n2117),
        .Q(n665) );
  AO22X1 U689 ( .IN1(n2119), .IN2(wr_data[10]), .IN3(\r[19][10] ), .IN4(n2117),
        .Q(n666) );
  AO22X1 U690 ( .IN1(n2119), .IN2(wr_data[11]), .IN3(\r[19][11] ), .IN4(n2117),
        .Q(n667) );
  AO22X1 U691 ( .IN1(n2119), .IN2(wr_data[12]), .IN3(\r[19][12] ), .IN4(n2117),
        .Q(n668) );
  AO22X1 U692 ( .IN1(n2119), .IN2(wr_data[13]), .IN3(\r[19][13] ), .IN4(n2117),
        .Q(n669) );
  AO22X1 U693 ( .IN1(n2119), .IN2(wr_data[14]), .IN3(\r[19][14] ), .IN4(n2117),
        .Q(n670) );
  AO22X1 U694 ( .IN1(n2119), .IN2(wr_data[15]), .IN3(\r[19][15] ), .IN4(n2117),
        .Q(n671) );
  AO22X1 U695 ( .IN1(n2119), .IN2(wr_data[16]), .IN3(\r[19][16] ), .IN4(n2117),
        .Q(n672) );
  AO22X1 U696 ( .IN1(n2119), .IN2(wr_data[17]), .IN3(\r[19][17] ), .IN4(n2117),
        .Q(n673) );
  AO22X1 U697 ( .IN1(n2119), .IN2(wr_data[18]), .IN3(\r[19][18] ), .IN4(n2117),
        .Q(n674) );
  AO22X1 U698 ( .IN1(n2119), .IN2(wr_data[19]), .IN3(\r[19][19] ), .IN4(n2117),
        .Q(n675) );
  AO22X1 U699 ( .IN1(n2119), .IN2(wr_data[20]), .IN3(\r[19][20] ), .IN4(n2116),
        .Q(n676) );
  AO22X1 U700 ( .IN1(n2119), .IN2(wr_data[21]), .IN3(\r[19][21] ), .IN4(n2116),
        .Q(n677) );
  AO22X1 U701 ( .IN1(n2119), .IN2(wr_data[22]), .IN3(\r[19][22] ), .IN4(n2116),
        .Q(n678) );
  AO22X1 U702 ( .IN1(n2120), .IN2(wr_data[23]), .IN3(\r[19][23] ), .IN4(n2116),
        .Q(n679) );
  AO22X1 U703 ( .IN1(n2120), .IN2(wr_data[24]), .IN3(\r[19][24] ), .IN4(n2116),
        .Q(n680) );
  AO22X1 U704 ( .IN1(n2120), .IN2(wr_data[25]), .IN3(\r[19][25] ), .IN4(n2116),
        .Q(n681) );
  AO22X1 U705 ( .IN1(n2120), .IN2(wr_data[26]), .IN3(\r[19][26] ), .IN4(n2116),
        .Q(n682) );
  AO22X1 U706 ( .IN1(n2120), .IN2(wr_data[27]), .IN3(\r[19][27] ), .IN4(n2116),
        .Q(n683) );
  AO22X1 U707 ( .IN1(n2120), .IN2(wr_data[28]), .IN3(\r[19][28] ), .IN4(n2116),
        .Q(n684) );
  AO22X1 U708 ( .IN1(n2120), .IN2(wr_data[29]), .IN3(\r[19][29] ), .IN4(n2116),
        .Q(n685) );
  AO22X1 U709 ( .IN1(n2120), .IN2(wr_data[30]), .IN3(\r[19][30] ), .IN4(n2116),
        .Q(n686) );
  AO22X1 U710 ( .IN1(n2120), .IN2(wr_data[31]), .IN3(\r[19][31] ), .IN4(n2116),
        .Q(n687) );
  AO22X1 U711 ( .IN1(n2113), .IN2(wr_data[0]), .IN3(\r[20][0] ), .IN4(n67),
        .Q(n688) );
  AO22X1 U712 ( .IN1(n2113), .IN2(wr_data[1]), .IN3(\r[20][1] ), .IN4(n67),
        .Q(n689) );
  AO22X1 U713 ( .IN1(n2113), .IN2(wr_data[2]), .IN3(\r[20][2] ), .IN4(n67),
        .Q(n690) );
  AO22X1 U714 ( .IN1(n2113), .IN2(wr_data[3]), .IN3(\r[20][3] ), .IN4(n67),
        .Q(n691) );
  AO22X1 U715 ( .IN1(n2113), .IN2(wr_data[4]), .IN3(\r[20][4] ), .IN4(n67),
        .Q(n692) );
  AO22X1 U716 ( .IN1(n2113), .IN2(wr_data[5]), .IN3(\r[20][5] ), .IN4(n67),
        .Q(n693) );
  AO22X1 U717 ( .IN1(n2113), .IN2(wr_data[6]), .IN3(\r[20][6] ), .IN4(n67),
        .Q(n694) );
  AO22X1 U718 ( .IN1(n2113), .IN2(wr_data[7]), .IN3(\r[20][7] ), .IN4(n67),
        .Q(n695) );
  AO22X1 U719 ( .IN1(n2113), .IN2(wr_data[8]), .IN3(\r[20][8] ), .IN4(n2112),
        .Q(n696) );
  AO22X1 U720 ( .IN1(n2113), .IN2(wr_data[9]), .IN3(\r[20][9] ), .IN4(n2112),
        .Q(n697) );
  AO22X1 U721 ( .IN1(n2114), .IN2(wr_data[10]), .IN3(\r[20][10] ), .IN4(n2112),
        .Q(n698) );
  AO22X1 U722 ( .IN1(n2114), .IN2(wr_data[11]), .IN3(\r[20][11] ), .IN4(n2112),
        .Q(n699) );
  AO22X1 U723 ( .IN1(n2114), .IN2(wr_data[12]), .IN3(\r[20][12] ), .IN4(n2112),
        .Q(n700) );
  AO22X1 U724 ( .IN1(n2114), .IN2(wr_data[13]), .IN3(\r[20][13] ), .IN4(n2112),
        .Q(n701) );
  AO22X1 U725 ( .IN1(n2114), .IN2(wr_data[14]), .IN3(\r[20][14] ), .IN4(n2112),
        .Q(n702) );
  AO22X1 U726 ( .IN1(n2114), .IN2(wr_data[15]), .IN3(\r[20][15] ), .IN4(n2112),
        .Q(n703) );
  AO22X1 U727 ( .IN1(n2114), .IN2(wr_data[16]), .IN3(\r[20][16] ), .IN4(n2112),
        .Q(n704) );
  AO22X1 U728 ( .IN1(n2114), .IN2(wr_data[17]), .IN3(\r[20][17] ), .IN4(n2112),
        .Q(n705) );
  AO22X1 U729 ( .IN1(n2114), .IN2(wr_data[18]), .IN3(\r[20][18] ), .IN4(n2112),
        .Q(n706) );
  AO22X1 U730 ( .IN1(n2114), .IN2(wr_data[19]), .IN3(\r[20][19] ), .IN4(n2112),
        .Q(n707) );
  AO22X1 U731 ( .IN1(n2114), .IN2(wr_data[20]), .IN3(\r[20][20] ), .IN4(n2111),
        .Q(n708) );
  AO22X1 U732 ( .IN1(n2114), .IN2(wr_data[21]), .IN3(\r[20][21] ), .IN4(n2111),
        .Q(n709) );
  AO22X1 U733 ( .IN1(n2114), .IN2(wr_data[22]), .IN3(\r[20][22] ), .IN4(n2111),
        .Q(n710) );
  AO22X1 U734 ( .IN1(n2115), .IN2(wr_data[23]), .IN3(\r[20][23] ), .IN4(n2111),
        .Q(n711) );
  AO22X1 U735 ( .IN1(n2115), .IN2(wr_data[24]), .IN3(\r[20][24] ), .IN4(n2111),
        .Q(n712) );
  AO22X1 U736 ( .IN1(n2115), .IN2(wr_data[25]), .IN3(\r[20][25] ), .IN4(n2111),
        .Q(n713) );
  AO22X1 U737 ( .IN1(n2115), .IN2(wr_data[26]), .IN3(\r[20][26] ), .IN4(n2111),
        .Q(n714) );
  AO22X1 U738 ( .IN1(n2115), .IN2(wr_data[27]), .IN3(\r[20][27] ), .IN4(n2111),
        .Q(n715) );
  AO22X1 U739 ( .IN1(n2115), .IN2(wr_data[28]), .IN3(\r[20][28] ), .IN4(n2111),
        .Q(n716) );
  AO22X1 U740 ( .IN1(n2115), .IN2(wr_data[29]), .IN3(\r[20][29] ), .IN4(n2111),
        .Q(n717) );
  AO22X1 U741 ( .IN1(n2115), .IN2(wr_data[30]), .IN3(\r[20][30] ), .IN4(n2111),
        .Q(n718) );
  AO22X1 U742 ( .IN1(n2115), .IN2(wr_data[31]), .IN3(\r[20][31] ), .IN4(n2111),
        .Q(n719) );
  AO22X1 U743 ( .IN1(n2108), .IN2(wr_data[0]), .IN3(\r[21][0] ), .IN4(n68),
        .Q(n720) );
  AO22X1 U744 ( .IN1(n2108), .IN2(wr_data[1]), .IN3(\r[21][1] ), .IN4(n68),
        .Q(n721) );
  AO22X1 U745 ( .IN1(n2108), .IN2(wr_data[2]), .IN3(\r[21][2] ), .IN4(n68),
        .Q(n722) );
  AO22X1 U746 ( .IN1(n2108), .IN2(wr_data[3]), .IN3(\r[21][3] ), .IN4(n68),
        .Q(n723) );
  AO22X1 U747 ( .IN1(n2108), .IN2(wr_data[4]), .IN3(\r[21][4] ), .IN4(n68),
        .Q(n724) );
  AO22X1 U748 ( .IN1(n2108), .IN2(wr_data[5]), .IN3(\r[21][5] ), .IN4(n68),
        .Q(n725) );
  AO22X1 U749 ( .IN1(n2108), .IN2(wr_data[6]), .IN3(\r[21][6] ), .IN4(n68),
        .Q(n726) );
  AO22X1 U750 ( .IN1(n2108), .IN2(wr_data[7]), .IN3(\r[21][7] ), .IN4(n68),
        .Q(n727) );
  AO22X1 U751 ( .IN1(n2108), .IN2(wr_data[8]), .IN3(\r[21][8] ), .IN4(n2107),
        .Q(n728) );
  AO22X1 U752 ( .IN1(n2108), .IN2(wr_data[9]), .IN3(\r[21][9] ), .IN4(n2107),
        .Q(n729) );
  AO22X1 U753 ( .IN1(n2109), .IN2(wr_data[10]), .IN3(\r[21][10] ), .IN4(n2107),
        .Q(n730) );
  AO22X1 U754 ( .IN1(n2109), .IN2(wr_data[11]), .IN3(\r[21][11] ), .IN4(n2107),
        .Q(n731) );
  AO22X1 U755 ( .IN1(n2109), .IN2(wr_data[12]), .IN3(\r[21][12] ), .IN4(n2107),
        .Q(n732) );
  AO22X1 U756 ( .IN1(n2109), .IN2(wr_data[13]), .IN3(\r[21][13] ), .IN4(n2107),
        .Q(n733) );
  AO22X1 U757 ( .IN1(n2109), .IN2(wr_data[14]), .IN3(\r[21][14] ), .IN4(n2107),
        .Q(n734) );
  AO22X1 U758 ( .IN1(n2109), .IN2(wr_data[15]), .IN3(\r[21][15] ), .IN4(n2107),
        .Q(n735) );
  AO22X1 U759 ( .IN1(n2109), .IN2(wr_data[16]), .IN3(\r[21][16] ), .IN4(n2107),
        .Q(n736) );
  AO22X1 U760 ( .IN1(n2109), .IN2(wr_data[17]), .IN3(\r[21][17] ), .IN4(n2107),
        .Q(n737) );
  AO22X1 U761 ( .IN1(n2109), .IN2(wr_data[18]), .IN3(\r[21][18] ), .IN4(n2107),
        .Q(n738) );
  AO22X1 U762 ( .IN1(n2109), .IN2(wr_data[19]), .IN3(\r[21][19] ), .IN4(n2107),
        .Q(n739) );
  AO22X1 U763 ( .IN1(n2109), .IN2(wr_data[20]), .IN3(\r[21][20] ), .IN4(n2106),
        .Q(n740) );
  AO22X1 U764 ( .IN1(n2109), .IN2(wr_data[21]), .IN3(\r[21][21] ), .IN4(n2106),
        .Q(n741) );
  AO22X1 U765 ( .IN1(n2109), .IN2(wr_data[22]), .IN3(\r[21][22] ), .IN4(n2106),
        .Q(n742) );
  AO22X1 U766 ( .IN1(n2110), .IN2(wr_data[23]), .IN3(\r[21][23] ), .IN4(n2106),
        .Q(n743) );
  AO22X1 U767 ( .IN1(n2110), .IN2(wr_data[24]), .IN3(\r[21][24] ), .IN4(n2106),
        .Q(n744) );
  AO22X1 U768 ( .IN1(n2110), .IN2(wr_data[25]), .IN3(\r[21][25] ), .IN4(n2106),
        .Q(n745) );
  AO22X1 U769 ( .IN1(n2110), .IN2(wr_data[26]), .IN3(\r[21][26] ), .IN4(n2106),
        .Q(n746) );
  AO22X1 U770 ( .IN1(n2110), .IN2(wr_data[27]), .IN3(\r[21][27] ), .IN4(n2106),
        .Q(n747) );
  AO22X1 U771 ( .IN1(n2110), .IN2(wr_data[28]), .IN3(\r[21][28] ), .IN4(n2106),
        .Q(n748) );
  AO22X1 U772 ( .IN1(n2110), .IN2(wr_data[29]), .IN3(\r[21][29] ), .IN4(n2106),
        .Q(n749) );
  AO22X1 U773 ( .IN1(n2110), .IN2(wr_data[30]), .IN3(\r[21][30] ), .IN4(n2106),
        .Q(n750) );
  AO22X1 U774 ( .IN1(n2110), .IN2(wr_data[31]), .IN3(\r[21][31] ), .IN4(n2106),
        .Q(n751) );
  AO22X1 U775 ( .IN1(n2103), .IN2(wr_data[0]), .IN3(\r[22][0] ), .IN4(n69),
        .Q(n752) );
  AO22X1 U776 ( .IN1(n2103), .IN2(wr_data[1]), .IN3(\r[22][1] ), .IN4(n69),
        .Q(n753) );
  AO22X1 U777 ( .IN1(n2103), .IN2(wr_data[2]), .IN3(\r[22][2] ), .IN4(n69),
        .Q(n754) );
  AO22X1 U778 ( .IN1(n2103), .IN2(wr_data[3]), .IN3(\r[22][3] ), .IN4(n69),
        .Q(n755) );
  AO22X1 U779 ( .IN1(n2103), .IN2(wr_data[4]), .IN3(\r[22][4] ), .IN4(n69),
        .Q(n756) );
  AO22X1 U780 ( .IN1(n2103), .IN2(wr_data[5]), .IN3(\r[22][5] ), .IN4(n69),
        .Q(n757) );
  AO22X1 U781 ( .IN1(n2103), .IN2(wr_data[6]), .IN3(\r[22][6] ), .IN4(n69),
        .Q(n758) );
  AO22X1 U782 ( .IN1(n2103), .IN2(wr_data[7]), .IN3(\r[22][7] ), .IN4(n69),
        .Q(n759) );
  AO22X1 U783 ( .IN1(n2103), .IN2(wr_data[8]), .IN3(\r[22][8] ), .IN4(n2102),
        .Q(n760) );
  AO22X1 U784 ( .IN1(n2103), .IN2(wr_data[9]), .IN3(\r[22][9] ), .IN4(n2102),
        .Q(n761) );
  AO22X1 U785 ( .IN1(n2104), .IN2(wr_data[10]), .IN3(\r[22][10] ), .IN4(n2102),
        .Q(n762) );
  AO22X1 U786 ( .IN1(n2104), .IN2(wr_data[11]), .IN3(\r[22][11] ), .IN4(n2102),
        .Q(n763) );
  AO22X1 U787 ( .IN1(n2104), .IN2(wr_data[12]), .IN3(\r[22][12] ), .IN4(n2102),
        .Q(n764) );
  AO22X1 U788 ( .IN1(n2104), .IN2(wr_data[13]), .IN3(\r[22][13] ), .IN4(n2102),
        .Q(n765) );
  AO22X1 U789 ( .IN1(n2104), .IN2(wr_data[14]), .IN3(\r[22][14] ), .IN4(n2102),
        .Q(n766) );
  AO22X1 U790 ( .IN1(n2104), .IN2(wr_data[15]), .IN3(\r[22][15] ), .IN4(n2102),
        .Q(n767) );
  AO22X1 U791 ( .IN1(n2104), .IN2(wr_data[16]), .IN3(\r[22][16] ), .IN4(n2102),
        .Q(n768) );
  AO22X1 U792 ( .IN1(n2104), .IN2(wr_data[17]), .IN3(\r[22][17] ), .IN4(n2102),
        .Q(n769) );
  AO22X1 U793 ( .IN1(n2104), .IN2(wr_data[18]), .IN3(\r[22][18] ), .IN4(n2102),
        .Q(n770) );
  AO22X1 U794 ( .IN1(n2104), .IN2(wr_data[19]), .IN3(\r[22][19] ), .IN4(n2102),
        .Q(n771) );
  AO22X1 U795 ( .IN1(n2104), .IN2(wr_data[20]), .IN3(\r[22][20] ), .IN4(n2101),
        .Q(n772) );
  AO22X1 U796 ( .IN1(n2104), .IN2(wr_data[21]), .IN3(\r[22][21] ), .IN4(n2101),
        .Q(n773) );
  AO22X1 U797 ( .IN1(n2104), .IN2(wr_data[22]), .IN3(\r[22][22] ), .IN4(n2101),
        .Q(n774) );
  AO22X1 U798 ( .IN1(n2105), .IN2(wr_data[23]), .IN3(\r[22][23] ), .IN4(n2101),
        .Q(n775) );
  AO22X1 U799 ( .IN1(n2105), .IN2(wr_data[24]), .IN3(\r[22][24] ), .IN4(n2101),
        .Q(n776) );
  AO22X1 U800 ( .IN1(n2105), .IN2(wr_data[25]), .IN3(\r[22][25] ), .IN4(n2101),
        .Q(n777) );
  AO22X1 U801 ( .IN1(n2105), .IN2(wr_data[26]), .IN3(\r[22][26] ), .IN4(n2101),
        .Q(n778) );
  AO22X1 U802 ( .IN1(n2105), .IN2(wr_data[27]), .IN3(\r[22][27] ), .IN4(n2101),
        .Q(n779) );
  AO22X1 U803 ( .IN1(n2105), .IN2(wr_data[28]), .IN3(\r[22][28] ), .IN4(n2101),
        .Q(n780) );
  AO22X1 U804 ( .IN1(n2105), .IN2(wr_data[29]), .IN3(\r[22][29] ), .IN4(n2101),
        .Q(n781) );
  AO22X1 U805 ( .IN1(n2105), .IN2(wr_data[30]), .IN3(\r[22][30] ), .IN4(n2101),
        .Q(n782) );
  AO22X1 U806 ( .IN1(n2105), .IN2(wr_data[31]), .IN3(\r[22][31] ), .IN4(n2101),
        .Q(n783) );
  AO22X1 U807 ( .IN1(n2098), .IN2(wr_data[0]), .IN3(\r[23][0] ), .IN4(n70),
        .Q(n784) );
  AO22X1 U808 ( .IN1(n2098), .IN2(wr_data[1]), .IN3(\r[23][1] ), .IN4(n70),
        .Q(n785) );
  AO22X1 U809 ( .IN1(n2098), .IN2(wr_data[2]), .IN3(\r[23][2] ), .IN4(n70),
        .Q(n786) );
  AO22X1 U810 ( .IN1(n2098), .IN2(wr_data[3]), .IN3(\r[23][3] ), .IN4(n70),
        .Q(n787) );
  AO22X1 U811 ( .IN1(n2098), .IN2(wr_data[4]), .IN3(\r[23][4] ), .IN4(n70),
        .Q(n788) );
  AO22X1 U812 ( .IN1(n2098), .IN2(wr_data[5]), .IN3(\r[23][5] ), .IN4(n70),
        .Q(n789) );
  AO22X1 U813 ( .IN1(n2098), .IN2(wr_data[6]), .IN3(\r[23][6] ), .IN4(n70),
        .Q(n790) );
  AO22X1 U814 ( .IN1(n2098), .IN2(wr_data[7]), .IN3(\r[23][7] ), .IN4(n70),
        .Q(n791) );
  AO22X1 U815 ( .IN1(n2098), .IN2(wr_data[8]), .IN3(\r[23][8] ), .IN4(n2097),
        .Q(n792) );
  AO22X1 U816 ( .IN1(n2098), .IN2(wr_data[9]), .IN3(\r[23][9] ), .IN4(n2097),
        .Q(n793) );
  AO22X1 U817 ( .IN1(n2099), .IN2(wr_data[10]), .IN3(\r[23][10] ), .IN4(n2097),
        .Q(n794) );
  AO22X1 U818 ( .IN1(n2099), .IN2(wr_data[11]), .IN3(\r[23][11] ), .IN4(n2097),
        .Q(n795) );
  AO22X1 U819 ( .IN1(n2099), .IN2(wr_data[12]), .IN3(\r[23][12] ), .IN4(n2097),
        .Q(n796) );
  AO22X1 U820 ( .IN1(n2099), .IN2(wr_data[13]), .IN3(\r[23][13] ), .IN4(n2097),
        .Q(n797) );
  AO22X1 U821 ( .IN1(n2099), .IN2(wr_data[14]), .IN3(\r[23][14] ), .IN4(n2097),
        .Q(n798) );
  AO22X1 U822 ( .IN1(n2099), .IN2(wr_data[15]), .IN3(\r[23][15] ), .IN4(n2097),
        .Q(n799) );
  AO22X1 U823 ( .IN1(n2099), .IN2(wr_data[16]), .IN3(\r[23][16] ), .IN4(n2097),
        .Q(n800) );
  AO22X1 U824 ( .IN1(n2099), .IN2(wr_data[17]), .IN3(\r[23][17] ), .IN4(n2097),
        .Q(n801) );
  AO22X1 U825 ( .IN1(n2099), .IN2(wr_data[18]), .IN3(\r[23][18] ), .IN4(n2097),
        .Q(n802) );
  AO22X1 U826 ( .IN1(n2099), .IN2(wr_data[19]), .IN3(\r[23][19] ), .IN4(n2097),
        .Q(n803) );
  AO22X1 U827 ( .IN1(n2099), .IN2(wr_data[20]), .IN3(\r[23][20] ), .IN4(n2096),
        .Q(n804) );
  AO22X1 U828 ( .IN1(n2099), .IN2(wr_data[21]), .IN3(\r[23][21] ), .IN4(n2096),
        .Q(n805) );
  AO22X1 U829 ( .IN1(n2099), .IN2(wr_data[22]), .IN3(\r[23][22] ), .IN4(n2096),
        .Q(n806) );
  AO22X1 U830 ( .IN1(n2100), .IN2(wr_data[23]), .IN3(\r[23][23] ), .IN4(n2096),
        .Q(n807) );
  AO22X1 U831 ( .IN1(n2100), .IN2(wr_data[24]), .IN3(\r[23][24] ), .IN4(n2096),
        .Q(n808) );
  AO22X1 U832 ( .IN1(n2100), .IN2(wr_data[25]), .IN3(\r[23][25] ), .IN4(n2096),
        .Q(n809) );
  AO22X1 U833 ( .IN1(n2100), .IN2(wr_data[26]), .IN3(\r[23][26] ), .IN4(n2096),
        .Q(n810) );
  AO22X1 U834 ( .IN1(n2100), .IN2(wr_data[27]), .IN3(\r[23][27] ), .IN4(n2096),
        .Q(n811) );
  AO22X1 U835 ( .IN1(n2100), .IN2(wr_data[28]), .IN3(\r[23][28] ), .IN4(n2096),
        .Q(n812) );
  AO22X1 U836 ( .IN1(n2100), .IN2(wr_data[29]), .IN3(\r[23][29] ), .IN4(n2096),
        .Q(n813) );
  AO22X1 U837 ( .IN1(n2100), .IN2(wr_data[30]), .IN3(\r[23][30] ), .IN4(n2096),
        .Q(n814) );
  AO22X1 U838 ( .IN1(n2100), .IN2(wr_data[31]), .IN3(\r[23][31] ), .IN4(n2096),
        .Q(n815) );
  AND3X1 U839 ( .IN1(wr_en), .IN2(n2300), .IN3(wr_addr[4]), .Q(n63) );
  AO22X1 U840 ( .IN1(n2093), .IN2(wr_data[0]), .IN3(\r[24][0] ), .IN4(n71),
        .Q(n816) );
  AO22X1 U841 ( .IN1(n2093), .IN2(wr_data[1]), .IN3(\r[24][1] ), .IN4(n71),
        .Q(n817) );
  AO22X1 U842 ( .IN1(n2093), .IN2(wr_data[2]), .IN3(\r[24][2] ), .IN4(n71),
        .Q(n818) );
  AO22X1 U843 ( .IN1(n2093), .IN2(wr_data[3]), .IN3(\r[24][3] ), .IN4(n71),
        .Q(n819) );
  AO22X1 U844 ( .IN1(n2093), .IN2(wr_data[4]), .IN3(\r[24][4] ), .IN4(n71),
        .Q(n820) );
  AO22X1 U845 ( .IN1(n2093), .IN2(wr_data[5]), .IN3(\r[24][5] ), .IN4(n71),
        .Q(n821) );
  AO22X1 U846 ( .IN1(n2093), .IN2(wr_data[6]), .IN3(\r[24][6] ), .IN4(n71),
        .Q(n822) );
  AO22X1 U847 ( .IN1(n2093), .IN2(wr_data[7]), .IN3(\r[24][7] ), .IN4(n71),
        .Q(n823) );
  AO22X1 U848 ( .IN1(n2093), .IN2(wr_data[8]), .IN3(\r[24][8] ), .IN4(n2092),
        .Q(n824) );
  AO22X1 U849 ( .IN1(n2093), .IN2(wr_data[9]), .IN3(\r[24][9] ), .IN4(n2092),
        .Q(n825) );
  AO22X1 U850 ( .IN1(n2094), .IN2(wr_data[10]), .IN3(\r[24][10] ), .IN4(n2092),
        .Q(n826) );
  AO22X1 U851 ( .IN1(n2094), .IN2(wr_data[11]), .IN3(\r[24][11] ), .IN4(n2092),
        .Q(n827) );
  AO22X1 U852 ( .IN1(n2094), .IN2(wr_data[12]), .IN3(\r[24][12] ), .IN4(n2092),
        .Q(n828) );
  AO22X1 U853 ( .IN1(n2094), .IN2(wr_data[13]), .IN3(\r[24][13] ), .IN4(n2092),
        .Q(n829) );
  AO22X1 U854 ( .IN1(n2094), .IN2(wr_data[14]), .IN3(\r[24][14] ), .IN4(n2092),
        .Q(n830) );
  AO22X1 U855 ( .IN1(n2094), .IN2(wr_data[15]), .IN3(\r[24][15] ), .IN4(n2092),
        .Q(n831) );
  AO22X1 U856 ( .IN1(n2094), .IN2(wr_data[16]), .IN3(\r[24][16] ), .IN4(n2092),
        .Q(n832) );
  AO22X1 U857 ( .IN1(n2094), .IN2(wr_data[17]), .IN3(\r[24][17] ), .IN4(n2092),
        .Q(n833) );
  AO22X1 U858 ( .IN1(n2094), .IN2(wr_data[18]), .IN3(\r[24][18] ), .IN4(n2092),
        .Q(n834) );
  AO22X1 U859 ( .IN1(n2094), .IN2(wr_data[19]), .IN3(\r[24][19] ), .IN4(n2092),
        .Q(n835) );
  AO22X1 U860 ( .IN1(n2094), .IN2(wr_data[20]), .IN3(\r[24][20] ), .IN4(n2091),
        .Q(n836) );
  AO22X1 U861 ( .IN1(n2094), .IN2(wr_data[21]), .IN3(\r[24][21] ), .IN4(n2091),
        .Q(n837) );
  AO22X1 U862 ( .IN1(n2094), .IN2(wr_data[22]), .IN3(\r[24][22] ), .IN4(n2091),
        .Q(n838) );
  AO22X1 U863 ( .IN1(n2095), .IN2(wr_data[23]), .IN3(\r[24][23] ), .IN4(n2091),
        .Q(n839) );
  AO22X1 U864 ( .IN1(n2095), .IN2(wr_data[24]), .IN3(\r[24][24] ), .IN4(n2091),
        .Q(n840) );
  AO22X1 U865 ( .IN1(n2095), .IN2(wr_data[25]), .IN3(\r[24][25] ), .IN4(n2091),
        .Q(n841) );
  AO22X1 U866 ( .IN1(n2095), .IN2(wr_data[26]), .IN3(\r[24][26] ), .IN4(n2091),
        .Q(n842) );
  AO22X1 U867 ( .IN1(n2095), .IN2(wr_data[27]), .IN3(\r[24][27] ), .IN4(n2091),
        .Q(n843) );
  AO22X1 U868 ( .IN1(n2095), .IN2(wr_data[28]), .IN3(\r[24][28] ), .IN4(n2091),
        .Q(n844) );
  AO22X1 U869 ( .IN1(n2095), .IN2(wr_data[29]), .IN3(\r[24][29] ), .IN4(n2091),
        .Q(n845) );
  AO22X1 U870 ( .IN1(n2095), .IN2(wr_data[30]), .IN3(\r[24][30] ), .IN4(n2091),
        .Q(n846) );
  AO22X1 U871 ( .IN1(n2095), .IN2(wr_data[31]), .IN3(\r[24][31] ), .IN4(n2091),
        .Q(n847) );
  AND3X1 U872 ( .IN1(n2302), .IN2(n2301), .IN3(n2303), .Q(n53) );
  AO22X1 U873 ( .IN1(n2088), .IN2(wr_data[0]), .IN3(\r[25][0] ), .IN4(n73),
        .Q(n848) );
  AO22X1 U874 ( .IN1(n2088), .IN2(wr_data[1]), .IN3(\r[25][1] ), .IN4(n73),
        .Q(n849) );
  AO22X1 U875 ( .IN1(n2088), .IN2(wr_data[2]), .IN3(\r[25][2] ), .IN4(n73),
        .Q(n850) );
  AO22X1 U876 ( .IN1(n2088), .IN2(wr_data[3]), .IN3(\r[25][3] ), .IN4(n73),
        .Q(n851) );
  AO22X1 U877 ( .IN1(n2088), .IN2(wr_data[4]), .IN3(\r[25][4] ), .IN4(n73),
        .Q(n852) );
  AO22X1 U878 ( .IN1(n2088), .IN2(wr_data[5]), .IN3(\r[25][5] ), .IN4(n73),
        .Q(n853) );
  AO22X1 U879 ( .IN1(n2088), .IN2(wr_data[6]), .IN3(\r[25][6] ), .IN4(n73),
        .Q(n854) );
  AO22X1 U880 ( .IN1(n2088), .IN2(wr_data[7]), .IN3(\r[25][7] ), .IN4(n73),
        .Q(n855) );
  AO22X1 U881 ( .IN1(n2088), .IN2(wr_data[8]), .IN3(\r[25][8] ), .IN4(n2087),
        .Q(n856) );
  AO22X1 U882 ( .IN1(n2088), .IN2(wr_data[9]), .IN3(\r[25][9] ), .IN4(n2087),
        .Q(n857) );
  AO22X1 U883 ( .IN1(n2089), .IN2(wr_data[10]), .IN3(\r[25][10] ), .IN4(n2087),
        .Q(n858) );
  AO22X1 U884 ( .IN1(n2089), .IN2(wr_data[11]), .IN3(\r[25][11] ), .IN4(n2087),
        .Q(n859) );
  AO22X1 U885 ( .IN1(n2089), .IN2(wr_data[12]), .IN3(\r[25][12] ), .IN4(n2087),
        .Q(n860) );
  AO22X1 U886 ( .IN1(n2089), .IN2(wr_data[13]), .IN3(\r[25][13] ), .IN4(n2087),
        .Q(n861) );
  AO22X1 U887 ( .IN1(n2089), .IN2(wr_data[14]), .IN3(\r[25][14] ), .IN4(n2087),
        .Q(n862) );
  AO22X1 U888 ( .IN1(n2089), .IN2(wr_data[15]), .IN3(\r[25][15] ), .IN4(n2087),
        .Q(n863) );
  AO22X1 U889 ( .IN1(n2089), .IN2(wr_data[16]), .IN3(\r[25][16] ), .IN4(n2087),
        .Q(n864) );
  AO22X1 U890 ( .IN1(n2089), .IN2(wr_data[17]), .IN3(\r[25][17] ), .IN4(n2087),
        .Q(n865) );
  AO22X1 U891 ( .IN1(n2089), .IN2(wr_data[18]), .IN3(\r[25][18] ), .IN4(n2087),
        .Q(n866) );
  AO22X1 U892 ( .IN1(n2089), .IN2(wr_data[19]), .IN3(\r[25][19] ), .IN4(n2087),
        .Q(n867) );
  AO22X1 U893 ( .IN1(n2089), .IN2(wr_data[20]), .IN3(\r[25][20] ), .IN4(n2086),
        .Q(n868) );
  AO22X1 U894 ( .IN1(n2089), .IN2(wr_data[21]), .IN3(\r[25][21] ), .IN4(n2086),
        .Q(n869) );
  AO22X1 U895 ( .IN1(n2089), .IN2(wr_data[22]), .IN3(\r[25][22] ), .IN4(n2086),
        .Q(n870) );
  AO22X1 U896 ( .IN1(n2090), .IN2(wr_data[23]), .IN3(\r[25][23] ), .IN4(n2086),
        .Q(n871) );
  AO22X1 U897 ( .IN1(n2090), .IN2(wr_data[24]), .IN3(\r[25][24] ), .IN4(n2086),
        .Q(n872) );
  AO22X1 U898 ( .IN1(n2090), .IN2(wr_data[25]), .IN3(\r[25][25] ), .IN4(n2086),
        .Q(n873) );
  AO22X1 U899 ( .IN1(n2090), .IN2(wr_data[26]), .IN3(\r[25][26] ), .IN4(n2086),
        .Q(n874) );
  AO22X1 U900 ( .IN1(n2090), .IN2(wr_data[27]), .IN3(\r[25][27] ), .IN4(n2086),
        .Q(n875) );
  AO22X1 U901 ( .IN1(n2090), .IN2(wr_data[28]), .IN3(\r[25][28] ), .IN4(n2086),
        .Q(n876) );
  AO22X1 U902 ( .IN1(n2090), .IN2(wr_data[29]), .IN3(\r[25][29] ), .IN4(n2086),
        .Q(n877) );
  AO22X1 U903 ( .IN1(n2090), .IN2(wr_data[30]), .IN3(\r[25][30] ), .IN4(n2086),
        .Q(n878) );
  AO22X1 U904 ( .IN1(n2090), .IN2(wr_data[31]), .IN3(\r[25][31] ), .IN4(n2086),
        .Q(n879) );
  AND3X1 U905 ( .IN1(n2302), .IN2(n2301), .IN3(wr_addr[0]), .Q(n38) );
  AO22X1 U906 ( .IN1(n2083), .IN2(wr_data[0]), .IN3(\r[26][0] ), .IN4(n74),
        .Q(n880) );
  AO22X1 U907 ( .IN1(n2083), .IN2(wr_data[1]), .IN3(\r[26][1] ), .IN4(n74),
        .Q(n881) );
  AO22X1 U908 ( .IN1(n2083), .IN2(wr_data[2]), .IN3(\r[26][2] ), .IN4(n74),
        .Q(n882) );
  AO22X1 U909 ( .IN1(n2083), .IN2(wr_data[3]), .IN3(\r[26][3] ), .IN4(n74),
        .Q(n883) );
  AO22X1 U910 ( .IN1(n2083), .IN2(wr_data[4]), .IN3(\r[26][4] ), .IN4(n74),
        .Q(n884) );
  AO22X1 U911 ( .IN1(n2083), .IN2(wr_data[5]), .IN3(\r[26][5] ), .IN4(n74),
        .Q(n885) );
  AO22X1 U912 ( .IN1(n2083), .IN2(wr_data[6]), .IN3(\r[26][6] ), .IN4(n74),
        .Q(n886) );
  AO22X1 U913 ( .IN1(n2083), .IN2(wr_data[7]), .IN3(\r[26][7] ), .IN4(n74),
        .Q(n887) );
  AO22X1 U914 ( .IN1(n2083), .IN2(wr_data[8]), .IN3(\r[26][8] ), .IN4(n2082),
        .Q(n888) );
  AO22X1 U915 ( .IN1(n2083), .IN2(wr_data[9]), .IN3(\r[26][9] ), .IN4(n2082),
        .Q(n889) );
  AO22X1 U916 ( .IN1(n2084), .IN2(wr_data[10]), .IN3(\r[26][10] ), .IN4(n2082),
        .Q(n890) );
  AO22X1 U917 ( .IN1(n2084), .IN2(wr_data[11]), .IN3(\r[26][11] ), .IN4(n2082),
        .Q(n891) );
  AO22X1 U918 ( .IN1(n2084), .IN2(wr_data[12]), .IN3(\r[26][12] ), .IN4(n2082),
        .Q(n892) );
  AO22X1 U919 ( .IN1(n2084), .IN2(wr_data[13]), .IN3(\r[26][13] ), .IN4(n2082),
        .Q(n893) );
  AO22X1 U920 ( .IN1(n2084), .IN2(wr_data[14]), .IN3(\r[26][14] ), .IN4(n2082),
        .Q(n894) );
  AO22X1 U921 ( .IN1(n2084), .IN2(wr_data[15]), .IN3(\r[26][15] ), .IN4(n2082),
        .Q(n895) );
  AO22X1 U922 ( .IN1(n2084), .IN2(wr_data[16]), .IN3(\r[26][16] ), .IN4(n2082),
        .Q(n896) );
  AO22X1 U923 ( .IN1(n2084), .IN2(wr_data[17]), .IN3(\r[26][17] ), .IN4(n2082),
        .Q(n897) );
  AO22X1 U924 ( .IN1(n2084), .IN2(wr_data[18]), .IN3(\r[26][18] ), .IN4(n2082),
        .Q(n898) );
  AO22X1 U925 ( .IN1(n2084), .IN2(wr_data[19]), .IN3(\r[26][19] ), .IN4(n2082),
        .Q(n899) );
  AO22X1 U926 ( .IN1(n2084), .IN2(wr_data[20]), .IN3(\r[26][20] ), .IN4(n2081),
        .Q(n900) );
  AO22X1 U927 ( .IN1(n2084), .IN2(wr_data[21]), .IN3(\r[26][21] ), .IN4(n2081),
        .Q(n901) );
  AO22X1 U928 ( .IN1(n2084), .IN2(wr_data[22]), .IN3(\r[26][22] ), .IN4(n2081),
        .Q(n902) );
  AO22X1 U929 ( .IN1(n2085), .IN2(wr_data[23]), .IN3(\r[26][23] ), .IN4(n2081),
        .Q(n903) );
  AO22X1 U930 ( .IN1(n2085), .IN2(wr_data[24]), .IN3(\r[26][24] ), .IN4(n2081),
        .Q(n904) );
  AO22X1 U931 ( .IN1(n2085), .IN2(wr_data[25]), .IN3(\r[26][25] ), .IN4(n2081),
        .Q(n905) );
  AO22X1 U932 ( .IN1(n2085), .IN2(wr_data[26]), .IN3(\r[26][26] ), .IN4(n2081),
        .Q(n906) );
  AO22X1 U933 ( .IN1(n2085), .IN2(wr_data[27]), .IN3(\r[26][27] ), .IN4(n2081),
        .Q(n907) );
  AO22X1 U934 ( .IN1(n2085), .IN2(wr_data[28]), .IN3(\r[26][28] ), .IN4(n2081),
        .Q(n908) );
  AO22X1 U935 ( .IN1(n2085), .IN2(wr_data[29]), .IN3(\r[26][29] ), .IN4(n2081),
        .Q(n909) );
  AO22X1 U936 ( .IN1(n2085), .IN2(wr_data[30]), .IN3(\r[26][30] ), .IN4(n2081),
        .Q(n910) );
  AO22X1 U937 ( .IN1(n2085), .IN2(wr_data[31]), .IN3(\r[26][31] ), .IN4(n2081),
        .Q(n911) );
  AND3X1 U938 ( .IN1(n2303), .IN2(n2301), .IN3(wr_addr[1]), .Q(n41) );
  AO22X1 U939 ( .IN1(n2078), .IN2(wr_data[0]), .IN3(\r[27][0] ), .IN4(n75),
        .Q(n912) );
  AO22X1 U940 ( .IN1(n2078), .IN2(wr_data[1]), .IN3(\r[27][1] ), .IN4(n75),
        .Q(n913) );
  AO22X1 U941 ( .IN1(n2078), .IN2(wr_data[2]), .IN3(\r[27][2] ), .IN4(n75),
        .Q(n914) );
  AO22X1 U942 ( .IN1(n2078), .IN2(wr_data[3]), .IN3(\r[27][3] ), .IN4(n75),
        .Q(n915) );
  AO22X1 U943 ( .IN1(n2078), .IN2(wr_data[4]), .IN3(\r[27][4] ), .IN4(n75),
        .Q(n916) );
  AO22X1 U944 ( .IN1(n2078), .IN2(wr_data[5]), .IN3(\r[27][5] ), .IN4(n75),
        .Q(n917) );
  AO22X1 U945 ( .IN1(n2078), .IN2(wr_data[6]), .IN3(\r[27][6] ), .IN4(n75),
        .Q(n918) );
  AO22X1 U946 ( .IN1(n2078), .IN2(wr_data[7]), .IN3(\r[27][7] ), .IN4(n75),
        .Q(n919) );
  AO22X1 U947 ( .IN1(n2078), .IN2(wr_data[8]), .IN3(\r[27][8] ), .IN4(n2077),
        .Q(n920) );
  AO22X1 U948 ( .IN1(n2078), .IN2(wr_data[9]), .IN3(\r[27][9] ), .IN4(n2077),
        .Q(n921) );
  AO22X1 U949 ( .IN1(n2079), .IN2(wr_data[10]), .IN3(\r[27][10] ), .IN4(n2077),
        .Q(n922) );
  AO22X1 U950 ( .IN1(n2079), .IN2(wr_data[11]), .IN3(\r[27][11] ), .IN4(n2077),
        .Q(n923) );
  AO22X1 U951 ( .IN1(n2079), .IN2(wr_data[12]), .IN3(\r[27][12] ), .IN4(n2077),
        .Q(n924) );
  AO22X1 U952 ( .IN1(n2079), .IN2(wr_data[13]), .IN3(\r[27][13] ), .IN4(n2077),
        .Q(n925) );
  AO22X1 U953 ( .IN1(n2079), .IN2(wr_data[14]), .IN3(\r[27][14] ), .IN4(n2077),
        .Q(n926) );
  AO22X1 U954 ( .IN1(n2079), .IN2(wr_data[15]), .IN3(\r[27][15] ), .IN4(n2077),
        .Q(n927) );
  AO22X1 U955 ( .IN1(n2079), .IN2(wr_data[16]), .IN3(\r[27][16] ), .IN4(n2077),
        .Q(n928) );
  AO22X1 U956 ( .IN1(n2079), .IN2(wr_data[17]), .IN3(\r[27][17] ), .IN4(n2077),
        .Q(n929) );
  AO22X1 U957 ( .IN1(n2079), .IN2(wr_data[18]), .IN3(\r[27][18] ), .IN4(n2077),
        .Q(n930) );
  AO22X1 U958 ( .IN1(n2079), .IN2(wr_data[19]), .IN3(\r[27][19] ), .IN4(n2077),
        .Q(n931) );
  AO22X1 U959 ( .IN1(n2079), .IN2(wr_data[20]), .IN3(\r[27][20] ), .IN4(n2076),
        .Q(n932) );
  AO22X1 U960 ( .IN1(n2079), .IN2(wr_data[21]), .IN3(\r[27][21] ), .IN4(n2076),
        .Q(n933) );
  AO22X1 U961 ( .IN1(n2079), .IN2(wr_data[22]), .IN3(\r[27][22] ), .IN4(n2076),
        .Q(n934) );
  AO22X1 U962 ( .IN1(n2080), .IN2(wr_data[23]), .IN3(\r[27][23] ), .IN4(n2076),
        .Q(n935) );
  AO22X1 U963 ( .IN1(n2080), .IN2(wr_data[24]), .IN3(\r[27][24] ), .IN4(n2076),
        .Q(n936) );
  AO22X1 U964 ( .IN1(n2080), .IN2(wr_data[25]), .IN3(\r[27][25] ), .IN4(n2076),
        .Q(n937) );
  AO22X1 U965 ( .IN1(n2080), .IN2(wr_data[26]), .IN3(\r[27][26] ), .IN4(n2076),
        .Q(n938) );
  AO22X1 U966 ( .IN1(n2080), .IN2(wr_data[27]), .IN3(\r[27][27] ), .IN4(n2076),
        .Q(n939) );
  AO22X1 U967 ( .IN1(n2080), .IN2(wr_data[28]), .IN3(\r[27][28] ), .IN4(n2076),
        .Q(n940) );
  AO22X1 U968 ( .IN1(n2080), .IN2(wr_data[29]), .IN3(\r[27][29] ), .IN4(n2076),
        .Q(n941) );
  AO22X1 U969 ( .IN1(n2080), .IN2(wr_data[30]), .IN3(\r[27][30] ), .IN4(n2076),
        .Q(n942) );
  AO22X1 U970 ( .IN1(n2080), .IN2(wr_data[31]), .IN3(\r[27][31] ), .IN4(n2076),
        .Q(n943) );
  AND3X1 U971 ( .IN1(wr_addr[0]), .IN2(n2301), .IN3(wr_addr[1]), .Q(n43) );
  AO22X1 U972 ( .IN1(n2073), .IN2(wr_data[0]), .IN3(\r[28][0] ), .IN4(n76),
        .Q(n944) );
  AO22X1 U973 ( .IN1(n2073), .IN2(wr_data[1]), .IN3(\r[28][1] ), .IN4(n76),
        .Q(n945) );
  AO22X1 U974 ( .IN1(n2073), .IN2(wr_data[2]), .IN3(\r[28][2] ), .IN4(n76),
        .Q(n946) );
  AO22X1 U975 ( .IN1(n2073), .IN2(wr_data[3]), .IN3(\r[28][3] ), .IN4(n76),
        .Q(n947) );
  AO22X1 U976 ( .IN1(n2073), .IN2(wr_data[4]), .IN3(\r[28][4] ), .IN4(n76),
        .Q(n948) );
  AO22X1 U977 ( .IN1(n2073), .IN2(wr_data[5]), .IN3(\r[28][5] ), .IN4(n76),
        .Q(n949) );
  AO22X1 U978 ( .IN1(n2073), .IN2(wr_data[6]), .IN3(\r[28][6] ), .IN4(n76),
        .Q(n950) );
  AO22X1 U979 ( .IN1(n2073), .IN2(wr_data[7]), .IN3(\r[28][7] ), .IN4(n76),
        .Q(n951) );
  AO22X1 U980 ( .IN1(n2073), .IN2(wr_data[8]), .IN3(\r[28][8] ), .IN4(n2072),
        .Q(n952) );
  AO22X1 U981 ( .IN1(n2073), .IN2(wr_data[9]), .IN3(\r[28][9] ), .IN4(n2072),
        .Q(n953) );
  AO22X1 U982 ( .IN1(n2074), .IN2(wr_data[10]), .IN3(\r[28][10] ), .IN4(n2072),
        .Q(n954) );
  AO22X1 U983 ( .IN1(n2074), .IN2(wr_data[11]), .IN3(\r[28][11] ), .IN4(n2072),
        .Q(n955) );
  AO22X1 U984 ( .IN1(n2074), .IN2(wr_data[12]), .IN3(\r[28][12] ), .IN4(n2072),
        .Q(n956) );
  AO22X1 U985 ( .IN1(n2074), .IN2(wr_data[13]), .IN3(\r[28][13] ), .IN4(n2072),
        .Q(n957) );
  AO22X1 U986 ( .IN1(n2074), .IN2(wr_data[14]), .IN3(\r[28][14] ), .IN4(n2072),
        .Q(n958) );
  AO22X1 U987 ( .IN1(n2074), .IN2(wr_data[15]), .IN3(\r[28][15] ), .IN4(n2072),
        .Q(n959) );
  AO22X1 U988 ( .IN1(n2074), .IN2(wr_data[16]), .IN3(\r[28][16] ), .IN4(n2072),
        .Q(n960) );
  AO22X1 U989 ( .IN1(n2074), .IN2(wr_data[17]), .IN3(\r[28][17] ), .IN4(n2072),
        .Q(n961) );
  AO22X1 U990 ( .IN1(n2074), .IN2(wr_data[18]), .IN3(\r[28][18] ), .IN4(n2072),
        .Q(n962) );
  AO22X1 U991 ( .IN1(n2074), .IN2(wr_data[19]), .IN3(\r[28][19] ), .IN4(n2072),
        .Q(n963) );
  AO22X1 U992 ( .IN1(n2074), .IN2(wr_data[20]), .IN3(\r[28][20] ), .IN4(n2071),
        .Q(n964) );
  AO22X1 U993 ( .IN1(n2074), .IN2(wr_data[21]), .IN3(\r[28][21] ), .IN4(n2071),
        .Q(n965) );
  AO22X1 U994 ( .IN1(n2074), .IN2(wr_data[22]), .IN3(\r[28][22] ), .IN4(n2071),
        .Q(n966) );
  AO22X1 U995 ( .IN1(n2075), .IN2(wr_data[23]), .IN3(\r[28][23] ), .IN4(n2071),
        .Q(n967) );
  AO22X1 U996 ( .IN1(n2075), .IN2(wr_data[24]), .IN3(\r[28][24] ), .IN4(n2071),
        .Q(n968) );
  AO22X1 U997 ( .IN1(n2075), .IN2(wr_data[25]), .IN3(\r[28][25] ), .IN4(n2071),
        .Q(n969) );
  AO22X1 U998 ( .IN1(n2075), .IN2(wr_data[26]), .IN3(\r[28][26] ), .IN4(n2071),
        .Q(n970) );
  AO22X1 U999 ( .IN1(n2075), .IN2(wr_data[27]), .IN3(\r[28][27] ), .IN4(n2071),
        .Q(n971) );
  AO22X1 U1000 ( .IN1(n2075), .IN2(wr_data[28]), .IN3(\r[28][28] ), .IN4(n2071), .Q(n972) );
  AO22X1 U1001 ( .IN1(n2075), .IN2(wr_data[29]), .IN3(\r[28][29] ), .IN4(n2071), .Q(n973) );
  AO22X1 U1002 ( .IN1(n2075), .IN2(wr_data[30]), .IN3(\r[28][30] ), .IN4(n2071), .Q(n974) );
  AO22X1 U1003 ( .IN1(n2075), .IN2(wr_data[31]), .IN3(\r[28][31] ), .IN4(n2071), .Q(n975) );
  AND3X1 U1004 ( .IN1(n2303), .IN2(n2302), .IN3(wr_addr[2]), .Q(n45) );
  AO22X1 U1005 ( .IN1(n2068), .IN2(wr_data[0]), .IN3(\r[29][0] ), .IN4(n77),
        .Q(n976) );
  AO22X1 U1006 ( .IN1(n2068), .IN2(wr_data[1]), .IN3(\r[29][1] ), .IN4(n77),
        .Q(n977) );
  AO22X1 U1007 ( .IN1(n2068), .IN2(wr_data[2]), .IN3(\r[29][2] ), .IN4(n77),
        .Q(n978) );
  AO22X1 U1008 ( .IN1(n2068), .IN2(wr_data[3]), .IN3(\r[29][3] ), .IN4(n77),
        .Q(n979) );
  AO22X1 U1009 ( .IN1(n2068), .IN2(wr_data[4]), .IN3(\r[29][4] ), .IN4(n77),
        .Q(n980) );
  AO22X1 U1010 ( .IN1(n2068), .IN2(wr_data[5]), .IN3(\r[29][5] ), .IN4(n77),
        .Q(n981) );
  AO22X1 U1011 ( .IN1(n2068), .IN2(wr_data[6]), .IN3(\r[29][6] ), .IN4(n77),
        .Q(n982) );
  AO22X1 U1012 ( .IN1(n2068), .IN2(wr_data[7]), .IN3(\r[29][7] ), .IN4(n77),
        .Q(n983) );
  AO22X1 U1013 ( .IN1(n2068), .IN2(wr_data[8]), .IN3(\r[29][8] ), .IN4(n2067),
        .Q(n984) );
  AO22X1 U1014 ( .IN1(n2068), .IN2(wr_data[9]), .IN3(\r[29][9] ), .IN4(n2067),
        .Q(n985) );
  AO22X1 U1015 ( .IN1(n2069), .IN2(wr_data[10]), .IN3(\r[29][10] ), .IN4(n2067), .Q(n986) );
  AO22X1 U1016 ( .IN1(n2069), .IN2(wr_data[11]), .IN3(\r[29][11] ), .IN4(n2067), .Q(n987) );
  AO22X1 U1017 ( .IN1(n2069), .IN2(wr_data[12]), .IN3(\r[29][12] ), .IN4(n2067), .Q(n988) );
  AO22X1 U1018 ( .IN1(n2069), .IN2(wr_data[13]), .IN3(\r[29][13] ), .IN4(n2067), .Q(n989) );
  AO22X1 U1019 ( .IN1(n2069), .IN2(wr_data[14]), .IN3(\r[29][14] ), .IN4(n2067), .Q(n990) );
  AO22X1 U1020 ( .IN1(n2069), .IN2(wr_data[15]), .IN3(\r[29][15] ), .IN4(n2067), .Q(n991) );
  AO22X1 U1021 ( .IN1(n2069), .IN2(wr_data[16]), .IN3(\r[29][16] ), .IN4(n2067), .Q(n992) );
  AO22X1 U1022 ( .IN1(n2069), .IN2(wr_data[17]), .IN3(\r[29][17] ), .IN4(n2067), .Q(n993) );
  AO22X1 U1023 ( .IN1(n2069), .IN2(wr_data[18]), .IN3(\r[29][18] ), .IN4(n2067), .Q(n994) );
  AO22X1 U1024 ( .IN1(n2069), .IN2(wr_data[19]), .IN3(\r[29][19] ), .IN4(n2067), .Q(n995) );
  AO22X1 U1025 ( .IN1(n2069), .IN2(wr_data[20]), .IN3(\r[29][20] ), .IN4(n2066), .Q(n996) );
  AO22X1 U1026 ( .IN1(n2069), .IN2(wr_data[21]), .IN3(\r[29][21] ), .IN4(n2066), .Q(n997) );
  AO22X1 U1027 ( .IN1(n2069), .IN2(wr_data[22]), .IN3(\r[29][22] ), .IN4(n2066), .Q(n998) );
  AO22X1 U1028 ( .IN1(n2070), .IN2(wr_data[23]), .IN3(\r[29][23] ), .IN4(n2066), .Q(n999) );
  AO22X1 U1029 ( .IN1(n2070), .IN2(wr_data[24]), .IN3(\r[29][24] ), .IN4(n2066), .Q(n1000) );
  AO22X1 U1030 ( .IN1(n2070), .IN2(wr_data[25]), .IN3(\r[29][25] ), .IN4(n2066), .Q(n1001) );
  AO22X1 U1031 ( .IN1(n2070), .IN2(wr_data[26]), .IN3(\r[29][26] ), .IN4(n2066), .Q(n1002) );
  AO22X1 U1032 ( .IN1(n2070), .IN2(wr_data[27]), .IN3(\r[29][27] ), .IN4(n2066), .Q(n1003) );
  AO22X1 U1033 ( .IN1(n2070), .IN2(wr_data[28]), .IN3(\r[29][28] ), .IN4(n2066), .Q(n1004) );
  AO22X1 U1034 ( .IN1(n2070), .IN2(wr_data[29]), .IN3(\r[29][29] ), .IN4(n2066), .Q(n1005) );
  AO22X1 U1035 ( .IN1(n2070), .IN2(wr_data[30]), .IN3(\r[29][30] ), .IN4(n2066), .Q(n1006) );
  AO22X1 U1036 ( .IN1(n2070), .IN2(wr_data[31]), .IN3(\r[29][31] ), .IN4(n2066), .Q(n1007) );
  AND3X1 U1037 ( .IN1(wr_addr[0]), .IN2(n2302), .IN3(wr_addr[2]), .Q(n47) );
  AO22X1 U1038 ( .IN1(n2063), .IN2(wr_data[0]), .IN3(\r[30][0] ), .IN4(n78),
        .Q(n1008) );
  AO22X1 U1039 ( .IN1(n2063), .IN2(wr_data[1]), .IN3(\r[30][1] ), .IN4(n78),
        .Q(n1009) );
  AO22X1 U1040 ( .IN1(n2063), .IN2(wr_data[2]), .IN3(\r[30][2] ), .IN4(n78),
        .Q(n1010) );
  AO22X1 U1041 ( .IN1(n2063), .IN2(wr_data[3]), .IN3(\r[30][3] ), .IN4(n78),
        .Q(n1011) );
  AO22X1 U1042 ( .IN1(n2063), .IN2(wr_data[4]), .IN3(\r[30][4] ), .IN4(n78),
        .Q(n1012) );
  AO22X1 U1043 ( .IN1(n2063), .IN2(wr_data[5]), .IN3(\r[30][5] ), .IN4(n78),
        .Q(n1013) );
  AO22X1 U1044 ( .IN1(n2063), .IN2(wr_data[6]), .IN3(\r[30][6] ), .IN4(n78),
        .Q(n1014) );
  AO22X1 U1045 ( .IN1(n2063), .IN2(wr_data[7]), .IN3(\r[30][7] ), .IN4(n78),
        .Q(n1015) );
  AO22X1 U1046 ( .IN1(n2063), .IN2(wr_data[8]), .IN3(\r[30][8] ), .IN4(n2062),
        .Q(n1016) );
  AO22X1 U1047 ( .IN1(n2063), .IN2(wr_data[9]), .IN3(\r[30][9] ), .IN4(n2062),
        .Q(n1017) );
  AO22X1 U1048 ( .IN1(n2064), .IN2(wr_data[10]), .IN3(\r[30][10] ), .IN4(n2062), .Q(n1018) );
  AO22X1 U1049 ( .IN1(n2064), .IN2(wr_data[11]), .IN3(\r[30][11] ), .IN4(n2062), .Q(n1019) );
  AO22X1 U1050 ( .IN1(n2064), .IN2(wr_data[12]), .IN3(\r[30][12] ), .IN4(n2062), .Q(n1020) );
  AO22X1 U1051 ( .IN1(n2064), .IN2(wr_data[13]), .IN3(\r[30][13] ), .IN4(n2062), .Q(n1021) );
  AO22X1 U1052 ( .IN1(n2064), .IN2(wr_data[14]), .IN3(\r[30][14] ), .IN4(n2062), .Q(n1022) );
  AO22X1 U1053 ( .IN1(n2064), .IN2(wr_data[15]), .IN3(\r[30][15] ), .IN4(n2062), .Q(n1023) );
  AO22X1 U1054 ( .IN1(n2064), .IN2(wr_data[16]), .IN3(\r[30][16] ), .IN4(n2062), .Q(n1024) );
  AO22X1 U1055 ( .IN1(n2064), .IN2(wr_data[17]), .IN3(\r[30][17] ), .IN4(n2062), .Q(n1025) );
  AO22X1 U1056 ( .IN1(n2064), .IN2(wr_data[18]), .IN3(\r[30][18] ), .IN4(n2062), .Q(n1026) );
  AO22X1 U1057 ( .IN1(n2064), .IN2(wr_data[19]), .IN3(\r[30][19] ), .IN4(n2062), .Q(n1027) );
  AO22X1 U1058 ( .IN1(n2064), .IN2(wr_data[20]), .IN3(\r[30][20] ), .IN4(n2061), .Q(n1028) );
  AO22X1 U1059 ( .IN1(n2064), .IN2(wr_data[21]), .IN3(\r[30][21] ), .IN4(n2061), .Q(n1029) );
  AO22X1 U1060 ( .IN1(n2064), .IN2(wr_data[22]), .IN3(\r[30][22] ), .IN4(n2061), .Q(n1030) );
  AO22X1 U1061 ( .IN1(n2065), .IN2(wr_data[23]), .IN3(\r[30][23] ), .IN4(n2061), .Q(n1031) );
  AO22X1 U1062 ( .IN1(n2065), .IN2(wr_data[24]), .IN3(\r[30][24] ), .IN4(n2061), .Q(n1032) );
  AO22X1 U1063 ( .IN1(n2065), .IN2(wr_data[25]), .IN3(\r[30][25] ), .IN4(n2061), .Q(n1033) );
  AO22X1 U1064 ( .IN1(n2065), .IN2(wr_data[26]), .IN3(\r[30][26] ), .IN4(n2061), .Q(n1034) );
  AO22X1 U1065 ( .IN1(n2065), .IN2(wr_data[27]), .IN3(\r[30][27] ), .IN4(n2061), .Q(n1035) );
  AO22X1 U1066 ( .IN1(n2065), .IN2(wr_data[28]), .IN3(\r[30][28] ), .IN4(n2061), .Q(n1036) );
  AO22X1 U1067 ( .IN1(n2065), .IN2(wr_data[29]), .IN3(\r[30][29] ), .IN4(n2061), .Q(n1037) );
  AO22X1 U1068 ( .IN1(n2065), .IN2(wr_data[30]), .IN3(\r[30][30] ), .IN4(n2061), .Q(n1038) );
  AO22X1 U1069 ( .IN1(n2065), .IN2(wr_data[31]), .IN3(\r[30][31] ), .IN4(n2061), .Q(n1039) );
  AND3X1 U1070 ( .IN1(wr_addr[1]), .IN2(n2303), .IN3(wr_addr[2]), .Q(n49) );
  AO22X1 U1071 ( .IN1(n2058), .IN2(wr_data[0]), .IN3(\r[31][0] ), .IN4(n79),
        .Q(n1040) );
  AO22X1 U1072 ( .IN1(n2058), .IN2(wr_data[1]), .IN3(\r[31][1] ), .IN4(n79),
        .Q(n1041) );
  AO22X1 U1073 ( .IN1(n2058), .IN2(wr_data[2]), .IN3(\r[31][2] ), .IN4(n79),
        .Q(n1042) );
  AO22X1 U1074 ( .IN1(n2058), .IN2(wr_data[3]), .IN3(\r[31][3] ), .IN4(n79),
        .Q(n1043) );
  AO22X1 U1075 ( .IN1(n2058), .IN2(wr_data[4]), .IN3(\r[31][4] ), .IN4(n79),
        .Q(n1044) );
  AO22X1 U1076 ( .IN1(n2058), .IN2(wr_data[5]), .IN3(\r[31][5] ), .IN4(n79),
        .Q(n1045) );
  AO22X1 U1077 ( .IN1(n2058), .IN2(wr_data[6]), .IN3(\r[31][6] ), .IN4(n79),
        .Q(n1046) );
  AO22X1 U1078 ( .IN1(n2058), .IN2(wr_data[7]), .IN3(\r[31][7] ), .IN4(n79),
        .Q(n1047) );
  AO22X1 U1079 ( .IN1(n2058), .IN2(wr_data[8]), .IN3(\r[31][8] ), .IN4(n2057),
        .Q(n1048) );
  AO22X1 U1080 ( .IN1(n2058), .IN2(wr_data[9]), .IN3(\r[31][9] ), .IN4(n2057),
        .Q(n1049) );
  AO22X1 U1081 ( .IN1(n2059), .IN2(wr_data[10]), .IN3(\r[31][10] ), .IN4(n2057), .Q(n1050) );
  AO22X1 U1082 ( .IN1(n2059), .IN2(wr_data[11]), .IN3(\r[31][11] ), .IN4(n2057), .Q(n1051) );
  AO22X1 U1083 ( .IN1(n2059), .IN2(wr_data[12]), .IN3(\r[31][12] ), .IN4(n2057), .Q(n1052) );
  AO22X1 U1084 ( .IN1(n2059), .IN2(wr_data[13]), .IN3(\r[31][13] ), .IN4(n2057), .Q(n1053) );
  AO22X1 U1085 ( .IN1(n2059), .IN2(wr_data[14]), .IN3(\r[31][14] ), .IN4(n2057), .Q(n1054) );
  AO22X1 U1086 ( .IN1(n2059), .IN2(wr_data[15]), .IN3(\r[31][15] ), .IN4(n2057), .Q(n1055) );
  AO22X1 U1087 ( .IN1(n2059), .IN2(wr_data[16]), .IN3(\r[31][16] ), .IN4(n2057), .Q(n1056) );
  AO22X1 U1088 ( .IN1(n2059), .IN2(wr_data[17]), .IN3(\r[31][17] ), .IN4(n2057), .Q(n1057) );
  AO22X1 U1089 ( .IN1(n2059), .IN2(wr_data[18]), .IN3(\r[31][18] ), .IN4(n2057), .Q(n1058) );
  AO22X1 U1090 ( .IN1(n2059), .IN2(wr_data[19]), .IN3(\r[31][19] ), .IN4(n2057), .Q(n1059) );
  AO22X1 U1091 ( .IN1(n2059), .IN2(wr_data[20]), .IN3(\r[31][20] ), .IN4(n2056), .Q(n1060) );
  AO22X1 U1092 ( .IN1(n2059), .IN2(wr_data[21]), .IN3(\r[31][21] ), .IN4(n2056), .Q(n1061) );
  AO22X1 U1093 ( .IN1(n2059), .IN2(wr_data[22]), .IN3(\r[31][22] ), .IN4(n2056), .Q(n1062) );
  AO22X1 U1094 ( .IN1(n2060), .IN2(wr_data[23]), .IN3(\r[31][23] ), .IN4(n2056), .Q(n1063) );
  AO22X1 U1095 ( .IN1(n2060), .IN2(wr_data[24]), .IN3(\r[31][24] ), .IN4(n2056), .Q(n1064) );
  AO22X1 U1096 ( .IN1(n2060), .IN2(wr_data[25]), .IN3(\r[31][25] ), .IN4(n2056), .Q(n1065) );
  AO22X1 U1097 ( .IN1(n2060), .IN2(wr_data[26]), .IN3(\r[31][26] ), .IN4(n2056), .Q(n1066) );
  AO22X1 U1098 ( .IN1(n2060), .IN2(wr_data[27]), .IN3(\r[31][27] ), .IN4(n2056), .Q(n1067) );
  AO22X1 U1099 ( .IN1(n2060), .IN2(wr_data[28]), .IN3(\r[31][28] ), .IN4(n2056), .Q(n1068) );
  AO22X1 U1100 ( .IN1(n2060), .IN2(wr_data[29]), .IN3(\r[31][29] ), .IN4(n2056), .Q(n1069) );
  AO22X1 U1101 ( .IN1(n2060), .IN2(wr_data[30]), .IN3(\r[31][30] ), .IN4(n2056), .Q(n1070) );
  AO22X1 U1102 ( .IN1(n2060), .IN2(wr_data[31]), .IN3(\r[31][31] ), .IN4(n2056), .Q(n1071) );
  AND3X1 U1103 ( .IN1(wr_addr[1]), .IN2(wr_addr[0]), .IN3(wr_addr[2]), .Q(n51)
         );
  AND3X1 U1104 ( .IN1(wr_addr[3]), .IN2(wr_en), .IN3(wr_addr[4]), .Q(n72) );
  INVX0 U1105 ( .INP(n55), .ZN(n2168) );
  INVX0 U1106 ( .INP(n56), .ZN(n2163) );
  INVX0 U1107 ( .INP(n57), .ZN(n2158) );
  INVX0 U1108 ( .INP(n58), .ZN(n2153) );
  INVX0 U1109 ( .INP(n59), .ZN(n2148) );
  INVX0 U1110 ( .INP(n60), .ZN(n2143) );
  INVX0 U1111 ( .INP(n61), .ZN(n2138) );
  INVX0 U1112 ( .INP(n62), .ZN(n2133) );
  INVX0 U1113 ( .INP(n64), .ZN(n2128) );
  INVX0 U1114 ( .INP(n65), .ZN(n2123) );
  INVX0 U1115 ( .INP(n66), .ZN(n2118) );
  INVX0 U1116 ( .INP(n67), .ZN(n2113) );
  INVX0 U1117 ( .INP(n68), .ZN(n2108) );
  INVX0 U1118 ( .INP(n69), .ZN(n2103) );
  INVX0 U1119 ( .INP(n70), .ZN(n2098) );
  INVX0 U1120 ( .INP(n71), .ZN(n2093) );
  INVX0 U1121 ( .INP(n73), .ZN(n2088) );
  INVX0 U1122 ( .INP(n74), .ZN(n2083) );
  INVX0 U1123 ( .INP(n75), .ZN(n2078) );
  INVX0 U1124 ( .INP(n76), .ZN(n2073) );
  INVX0 U1125 ( .INP(n77), .ZN(n2068) );
  INVX0 U1126 ( .INP(n78), .ZN(n2063) );
  INVX0 U1127 ( .INP(n79), .ZN(n2058) );
  INVX0 U1128 ( .INP(n52), .ZN(n2173) );
  INVX0 U1129 ( .INP(n37), .ZN(n2208) );
  INVX0 U1130 ( .INP(n40), .ZN(n2203) );
  INVX0 U1131 ( .INP(n42), .ZN(n2198) );
  INVX0 U1132 ( .INP(n44), .ZN(n2193) );
  INVX0 U1133 ( .INP(n46), .ZN(n2188) );
  INVX0 U1134 ( .INP(n48), .ZN(n2183) );
  INVX0 U1135 ( .INP(n50), .ZN(n2178) );
  INVX0 U1136 ( .INP(N17), .ZN(n2035) );
  INVX0 U1137 ( .INP(N12), .ZN(n1543) );
  INVX0 U1138 ( .INP(N16), .ZN(n2013) );
  INVX0 U1139 ( .INP(N11), .ZN(n1521) );
  INVX0 U1140 ( .INP(N16), .ZN(n2012) );
  INVX0 U1141 ( .INP(N11), .ZN(n1520) );
  INVX0 U1142 ( .INP(N18), .ZN(n2051) );
  INVX0 U1143 ( .INP(N13), .ZN(n1559) );
  INVX0 U1144 ( .INP(n2173), .ZN(n2172) );
  INVX0 U1145 ( .INP(n2173), .ZN(n2171) );
  INVX0 U1146 ( .INP(n2203), .ZN(n2202) );
  INVX0 U1147 ( .INP(n2203), .ZN(n2201) );
  INVX0 U1148 ( .INP(n2198), .ZN(n2197) );
  INVX0 U1149 ( .INP(n2198), .ZN(n2196) );
  INVX0 U1150 ( .INP(n2193), .ZN(n2192) );
  INVX0 U1151 ( .INP(n2193), .ZN(n2191) );
  INVX0 U1152 ( .INP(n2188), .ZN(n2187) );
  INVX0 U1153 ( .INP(n2188), .ZN(n2186) );
  INVX0 U1154 ( .INP(n2183), .ZN(n2182) );
  INVX0 U1155 ( .INP(n2183), .ZN(n2181) );
  INVX0 U1156 ( .INP(n2178), .ZN(n2177) );
  INVX0 U1157 ( .INP(n2178), .ZN(n2176) );
  INVX0 U1158 ( .INP(n2208), .ZN(n2207) );
  INVX0 U1159 ( .INP(n2208), .ZN(n2206) );
  INVX0 U1160 ( .INP(n2133), .ZN(n2132) );
  INVX0 U1161 ( .INP(n2133), .ZN(n2131) );
  INVX0 U1162 ( .INP(n2128), .ZN(n2127) );
  INVX0 U1163 ( .INP(n2128), .ZN(n2126) );
  INVX0 U1164 ( .INP(n2123), .ZN(n2122) );
  INVX0 U1165 ( .INP(n2123), .ZN(n2121) );
  INVX0 U1166 ( .INP(n2118), .ZN(n2117) );
  INVX0 U1167 ( .INP(n2118), .ZN(n2116) );
  INVX0 U1168 ( .INP(n2113), .ZN(n2112) );
  INVX0 U1169 ( .INP(n2113), .ZN(n2111) );
  INVX0 U1170 ( .INP(n2108), .ZN(n2107) );
  INVX0 U1171 ( .INP(n2108), .ZN(n2106) );
  INVX0 U1172 ( .INP(n2103), .ZN(n2102) );
  INVX0 U1173 ( .INP(n2103), .ZN(n2101) );
  INVX0 U1174 ( .INP(n2098), .ZN(n2097) );
  INVX0 U1175 ( .INP(n2098), .ZN(n2096) );
  INVX0 U1176 ( .INP(n2093), .ZN(n2092) );
  INVX0 U1177 ( .INP(n2093), .ZN(n2091) );
  INVX0 U1178 ( .INP(n2088), .ZN(n2087) );
  INVX0 U1179 ( .INP(n2088), .ZN(n2086) );
  INVX0 U1180 ( .INP(n2083), .ZN(n2082) );
  INVX0 U1181 ( .INP(n2083), .ZN(n2081) );
  INVX0 U1182 ( .INP(n2078), .ZN(n2077) );
  INVX0 U1183 ( .INP(n2078), .ZN(n2076) );
  INVX0 U1184 ( .INP(n2073), .ZN(n2072) );
  INVX0 U1185 ( .INP(n2073), .ZN(n2071) );
  INVX0 U1186 ( .INP(n2068), .ZN(n2067) );
  INVX0 U1187 ( .INP(n2068), .ZN(n2066) );
  INVX0 U1188 ( .INP(n2063), .ZN(n2062) );
  INVX0 U1189 ( .INP(n2063), .ZN(n2061) );
  INVX0 U1190 ( .INP(n2058), .ZN(n2057) );
  INVX0 U1191 ( .INP(n2058), .ZN(n2056) );
  INVX0 U1192 ( .INP(n2168), .ZN(n2167) );
  INVX0 U1193 ( .INP(n2168), .ZN(n2166) );
  INVX0 U1194 ( .INP(n2163), .ZN(n2162) );
  INVX0 U1195 ( .INP(n2163), .ZN(n2161) );
  INVX0 U1196 ( .INP(n2158), .ZN(n2157) );
  INVX0 U1197 ( .INP(n2158), .ZN(n2156) );
  INVX0 U1198 ( .INP(n2153), .ZN(n2152) );
  INVX0 U1199 ( .INP(n2153), .ZN(n2151) );
  INVX0 U1200 ( .INP(n2148), .ZN(n2147) );
  INVX0 U1201 ( .INP(n2148), .ZN(n2146) );
  INVX0 U1202 ( .INP(n2143), .ZN(n2142) );
  INVX0 U1203 ( .INP(n2143), .ZN(n2141) );
  INVX0 U1204 ( .INP(n2138), .ZN(n2137) );
  INVX0 U1205 ( .INP(n2138), .ZN(n2136) );
  INVX0 U1206 ( .INP(n52), .ZN(n2174) );
  INVX0 U1207 ( .INP(n40), .ZN(n2204) );
  INVX0 U1208 ( .INP(n42), .ZN(n2199) );
  INVX0 U1209 ( .INP(n44), .ZN(n2194) );
  INVX0 U1210 ( .INP(n46), .ZN(n2189) );
  INVX0 U1211 ( .INP(n48), .ZN(n2184) );
  INVX0 U1212 ( .INP(n50), .ZN(n2179) );
  INVX0 U1213 ( .INP(n37), .ZN(n2209) );
  INVX0 U1214 ( .INP(n62), .ZN(n2134) );
  INVX0 U1215 ( .INP(n64), .ZN(n2129) );
  INVX0 U1216 ( .INP(n65), .ZN(n2124) );
  INVX0 U1217 ( .INP(n66), .ZN(n2119) );
  INVX0 U1218 ( .INP(n67), .ZN(n2114) );
  INVX0 U1219 ( .INP(n68), .ZN(n2109) );
  INVX0 U1220 ( .INP(n69), .ZN(n2104) );
  INVX0 U1221 ( .INP(n70), .ZN(n2099) );
  INVX0 U1222 ( .INP(n71), .ZN(n2094) );
  INVX0 U1223 ( .INP(n73), .ZN(n2089) );
  INVX0 U1224 ( .INP(n74), .ZN(n2084) );
  INVX0 U1225 ( .INP(n75), .ZN(n2079) );
  INVX0 U1226 ( .INP(n76), .ZN(n2074) );
  INVX0 U1227 ( .INP(n77), .ZN(n2069) );
  INVX0 U1228 ( .INP(n78), .ZN(n2064) );
  INVX0 U1229 ( .INP(n79), .ZN(n2059) );
  INVX0 U1230 ( .INP(n55), .ZN(n2169) );
  INVX0 U1231 ( .INP(n56), .ZN(n2164) );
  INVX0 U1232 ( .INP(n57), .ZN(n2159) );
  INVX0 U1233 ( .INP(n58), .ZN(n2154) );
  INVX0 U1234 ( .INP(n59), .ZN(n2149) );
  INVX0 U1235 ( .INP(n60), .ZN(n2144) );
  INVX0 U1236 ( .INP(n61), .ZN(n2139) );
  INVX0 U1237 ( .INP(n52), .ZN(n2175) );
  INVX0 U1238 ( .INP(n40), .ZN(n2205) );
  INVX0 U1239 ( .INP(n42), .ZN(n2200) );
  INVX0 U1240 ( .INP(n44), .ZN(n2195) );
  INVX0 U1241 ( .INP(n46), .ZN(n2190) );
  INVX0 U1242 ( .INP(n48), .ZN(n2185) );
  INVX0 U1243 ( .INP(n50), .ZN(n2180) );
  INVX0 U1244 ( .INP(n37), .ZN(n2210) );
  INVX0 U1245 ( .INP(n62), .ZN(n2135) );
  INVX0 U1246 ( .INP(n64), .ZN(n2130) );
  INVX0 U1247 ( .INP(n65), .ZN(n2125) );
  INVX0 U1248 ( .INP(n66), .ZN(n2120) );
  INVX0 U1249 ( .INP(n67), .ZN(n2115) );
  INVX0 U1250 ( .INP(n68), .ZN(n2110) );
  INVX0 U1251 ( .INP(n69), .ZN(n2105) );
  INVX0 U1252 ( .INP(n70), .ZN(n2100) );
  INVX0 U1253 ( .INP(n71), .ZN(n2095) );
  INVX0 U1254 ( .INP(n73), .ZN(n2090) );
  INVX0 U1255 ( .INP(n74), .ZN(n2085) );
  INVX0 U1256 ( .INP(n75), .ZN(n2080) );
  INVX0 U1257 ( .INP(n76), .ZN(n2075) );
  INVX0 U1258 ( .INP(n77), .ZN(n2070) );
  INVX0 U1259 ( .INP(n78), .ZN(n2065) );
  INVX0 U1260 ( .INP(n79), .ZN(n2060) );
  INVX0 U1261 ( .INP(n55), .ZN(n2170) );
  INVX0 U1262 ( .INP(n56), .ZN(n2165) );
  INVX0 U1263 ( .INP(n57), .ZN(n2160) );
  INVX0 U1264 ( .INP(n58), .ZN(n2155) );
  INVX0 U1265 ( .INP(n59), .ZN(n2150) );
  INVX0 U1266 ( .INP(n60), .ZN(n2145) );
  INVX0 U1267 ( .INP(n61), .ZN(n2140) );
  INVX0 U1268 ( .INP(n2035), .ZN(n2049) );
  INVX0 U1269 ( .INP(n1543), .ZN(n1557) );
  INVX0 U1270 ( .INP(n2035), .ZN(n2050) );
  INVX0 U1271 ( .INP(n1543), .ZN(n1558) );
  INVX0 U1272 ( .INP(n2035), .ZN(n2044) );
  INVX0 U1273 ( .INP(n2035), .ZN(n2045) );
  INVX0 U1274 ( .INP(n2035), .ZN(n2047) );
  INVX0 U1275 ( .INP(n2035), .ZN(n2048) );
  INVX0 U1276 ( .INP(n2035), .ZN(n2046) );
  INVX0 U1277 ( .INP(n2035), .ZN(n2040) );
  INVX0 U1278 ( .INP(n2035), .ZN(n2041) );
  INVX0 U1279 ( .INP(n2035), .ZN(n2042) );
  INVX0 U1280 ( .INP(n2035), .ZN(n2043) );
  INVX0 U1281 ( .INP(n1543), .ZN(n1552) );
  INVX0 U1282 ( .INP(n1543), .ZN(n1553) );
  INVX0 U1283 ( .INP(n1543), .ZN(n1555) );
  INVX0 U1284 ( .INP(n1543), .ZN(n1556) );
  INVX0 U1285 ( .INP(n1543), .ZN(n1554) );
  INVX0 U1286 ( .INP(n1543), .ZN(n1548) );
  INVX0 U1287 ( .INP(n1543), .ZN(n1549) );
  INVX0 U1288 ( .INP(n1543), .ZN(n1550) );
  INVX0 U1289 ( .INP(n1543), .ZN(n1551) );
  INVX0 U1290 ( .INP(n2013), .ZN(n2016) );
  INVX0 U1291 ( .INP(n1521), .ZN(n1524) );
  INVX0 U1292 ( .INP(n2013), .ZN(n2015) );
  INVX0 U1293 ( .INP(n1521), .ZN(n1523) );
  INVX0 U1294 ( .INP(n2013), .ZN(n2017) );
  INVX0 U1295 ( .INP(n1521), .ZN(n1525) );
  INVX0 U1296 ( .INP(n2013), .ZN(n2024) );
  INVX0 U1297 ( .INP(n2013), .ZN(n2018) );
  INVX0 U1298 ( .INP(n2013), .ZN(n2019) );
  INVX0 U1299 ( .INP(n2013), .ZN(n2020) );
  INVX0 U1300 ( .INP(n2013), .ZN(n2021) );
  INVX0 U1301 ( .INP(n2013), .ZN(n2022) );
  INVX0 U1302 ( .INP(n2013), .ZN(n2023) );
  INVX0 U1303 ( .INP(n1521), .ZN(n1532) );
  INVX0 U1304 ( .INP(n1521), .ZN(n1526) );
  INVX0 U1305 ( .INP(n1521), .ZN(n1527) );
  INVX0 U1306 ( .INP(n1521), .ZN(n1528) );
  INVX0 U1307 ( .INP(n1521), .ZN(n1529) );
  INVX0 U1308 ( .INP(n1521), .ZN(n1530) );
  INVX0 U1309 ( .INP(n1521), .ZN(n1531) );
  INVX0 U1310 ( .INP(n2013), .ZN(n2014) );
  INVX0 U1311 ( .INP(n1521), .ZN(n1522) );
  INVX0 U1312 ( .INP(n2012), .ZN(n2025) );
  INVX0 U1313 ( .INP(n2012), .ZN(n2026) );
  INVX0 U1314 ( .INP(n2012), .ZN(n2027) );
  INVX0 U1315 ( .INP(n2012), .ZN(n2028) );
  INVX0 U1316 ( .INP(n2012), .ZN(n2030) );
  INVX0 U1317 ( .INP(n2012), .ZN(n2031) );
  INVX0 U1318 ( .INP(n2012), .ZN(n2032) );
  INVX0 U1319 ( .INP(n2012), .ZN(n2033) );
  INVX0 U1320 ( .INP(n2012), .ZN(n2029) );
  INVX0 U1321 ( .INP(n2012), .ZN(n2034) );
  INVX0 U1322 ( .INP(n1520), .ZN(n1533) );
  INVX0 U1323 ( .INP(n1520), .ZN(n1534) );
  INVX0 U1324 ( .INP(n1520), .ZN(n1535) );
  INVX0 U1325 ( .INP(n1520), .ZN(n1536) );
  INVX0 U1326 ( .INP(n1520), .ZN(n1538) );
  INVX0 U1327 ( .INP(n1520), .ZN(n1539) );
  INVX0 U1328 ( .INP(n1520), .ZN(n1540) );
  INVX0 U1329 ( .INP(n1520), .ZN(n1541) );
  INVX0 U1330 ( .INP(n1520), .ZN(n1537) );
  INVX0 U1331 ( .INP(n1520), .ZN(n1542) );
  INVX0 U1332 ( .INP(n2051), .ZN(n2055) );
  INVX0 U1333 ( .INP(n2051), .ZN(n2054) );
  INVX0 U1334 ( .INP(n2051), .ZN(n2053) );
  INVX0 U1335 ( .INP(n1559), .ZN(n1563) );
  INVX0 U1336 ( .INP(n1559), .ZN(n1562) );
  INVX0 U1337 ( .INP(n1559), .ZN(n1561) );
  INVX0 U1338 ( .INP(n2051), .ZN(n2052) );
  INVX0 U1339 ( .INP(n1559), .ZN(n1560) );
  INVX0 U1340 ( .INP(n2037), .ZN(n2039) );
  INVX0 U1341 ( .INP(n1545), .ZN(n1547) );
  INVX0 U1342 ( .INP(n2036), .ZN(n2038) );
  INVX0 U1343 ( .INP(n1544), .ZN(n1546) );
  NAND2X1 U1344 ( .IN1(n53), .IN2(n54), .QN(n52) );
  NAND2X1 U1345 ( .IN1(n38), .IN2(n39), .QN(n37) );
  NAND2X1 U1346 ( .IN1(n41), .IN2(n39), .QN(n40) );
  NAND2X1 U1347 ( .IN1(n43), .IN2(n39), .QN(n42) );
  NAND2X1 U1348 ( .IN1(n45), .IN2(n39), .QN(n44) );
  NAND2X1 U1349 ( .IN1(n47), .IN2(n39), .QN(n46) );
  NAND2X1 U1350 ( .IN1(n49), .IN2(n39), .QN(n48) );
  NAND2X1 U1351 ( .IN1(n51), .IN2(n39), .QN(n50) );
  NAND2X1 U1352 ( .IN1(n63), .IN2(n53), .QN(n62) );
  NAND2X1 U1353 ( .IN1(n63), .IN2(n38), .QN(n64) );
  NAND2X1 U1354 ( .IN1(n63), .IN2(n41), .QN(n65) );
  NAND2X1 U1355 ( .IN1(n63), .IN2(n43), .QN(n66) );
  NAND2X1 U1356 ( .IN1(n63), .IN2(n45), .QN(n67) );
  NAND2X1 U1357 ( .IN1(n63), .IN2(n47), .QN(n68) );
  NAND2X1 U1358 ( .IN1(n63), .IN2(n49), .QN(n69) );
  NAND2X1 U1359 ( .IN1(n63), .IN2(n51), .QN(n70) );
  NAND2X1 U1360 ( .IN1(n72), .IN2(n53), .QN(n71) );
  NAND2X1 U1361 ( .IN1(n72), .IN2(n38), .QN(n73) );
  NAND2X1 U1362 ( .IN1(n72), .IN2(n41), .QN(n74) );
  NAND2X1 U1363 ( .IN1(n72), .IN2(n43), .QN(n75) );
  NAND2X1 U1364 ( .IN1(n72), .IN2(n45), .QN(n76) );
  NAND2X1 U1365 ( .IN1(n72), .IN2(n47), .QN(n77) );
  NAND2X1 U1366 ( .IN1(n72), .IN2(n49), .QN(n78) );
  NAND2X1 U1367 ( .IN1(n72), .IN2(n51), .QN(n79) );
  NAND2X1 U1368 ( .IN1(n54), .IN2(n38), .QN(n55) );
  NAND2X1 U1369 ( .IN1(n54), .IN2(n41), .QN(n56) );
  NAND2X1 U1370 ( .IN1(n54), .IN2(n43), .QN(n57) );
  NAND2X1 U1371 ( .IN1(n54), .IN2(n45), .QN(n58) );
  NAND2X1 U1372 ( .IN1(n54), .IN2(n47), .QN(n59) );
  NAND2X1 U1373 ( .IN1(n54), .IN2(n49), .QN(n60) );
  NAND2X1 U1374 ( .IN1(n54), .IN2(n51), .QN(n61) );
  INVX0 U1375 ( .INP(n2293), .ZN(n2221) );
  INVX0 U1376 ( .INP(n2294), .ZN(n2220) );
  INVX0 U1377 ( .INP(n2295), .ZN(n2219) );
  INVX0 U1378 ( .INP(n2296), .ZN(n2218) );
  INVX0 U1379 ( .INP(n2297), .ZN(n2217) );
  INVX0 U1380 ( .INP(n2298), .ZN(n2216) );
  INVX0 U1381 ( .INP(n2293), .ZN(n2215) );
  INVX0 U1382 ( .INP(n2294), .ZN(n2214) );
  INVX0 U1383 ( .INP(n2295), .ZN(n2213) );
  INVX0 U1384 ( .INP(n2296), .ZN(n2212) );
  INVX0 U1385 ( .INP(n2297), .ZN(n2211) );
  INVX0 U1386 ( .INP(n2293), .ZN(n2292) );
  INVX0 U1387 ( .INP(n2293), .ZN(n2291) );
  INVX0 U1388 ( .INP(n2293), .ZN(n2290) );
  INVX0 U1389 ( .INP(n2293), .ZN(n2289) );
  INVX0 U1390 ( .INP(n2293), .ZN(n2288) );
  INVX0 U1391 ( .INP(n2293), .ZN(n2287) );
  INVX0 U1392 ( .INP(n2293), .ZN(n2286) );
  INVX0 U1393 ( .INP(n2293), .ZN(n2285) );
  INVX0 U1394 ( .INP(n2293), .ZN(n2284) );
  INVX0 U1395 ( .INP(n2293), .ZN(n2283) );
  INVX0 U1396 ( .INP(n2293), .ZN(n2282) );
  INVX0 U1397 ( .INP(n2294), .ZN(n2281) );
  INVX0 U1398 ( .INP(n2294), .ZN(n2280) );
  INVX0 U1399 ( .INP(n2294), .ZN(n2279) );
  INVX0 U1400 ( .INP(n2294), .ZN(n2278) );
  INVX0 U1401 ( .INP(n2294), .ZN(n2277) );
  INVX0 U1402 ( .INP(n2294), .ZN(n2276) );
  INVX0 U1403 ( .INP(n2294), .ZN(n2275) );
  INVX0 U1404 ( .INP(n2294), .ZN(n2274) );
  INVX0 U1405 ( .INP(n2294), .ZN(n2273) );
  INVX0 U1406 ( .INP(n2294), .ZN(n2272) );
  INVX0 U1407 ( .INP(n2294), .ZN(n2271) );
  INVX0 U1408 ( .INP(n2294), .ZN(n2270) );
  INVX0 U1409 ( .INP(n2295), .ZN(n2269) );
  INVX0 U1410 ( .INP(n2295), .ZN(n2268) );
  INVX0 U1411 ( .INP(n2295), .ZN(n2267) );
  INVX0 U1412 ( .INP(n2295), .ZN(n2266) );
  INVX0 U1413 ( .INP(n2295), .ZN(n2265) );
  INVX0 U1414 ( .INP(n2295), .ZN(n2264) );
  INVX0 U1415 ( .INP(n2295), .ZN(n2263) );
  INVX0 U1416 ( .INP(n2295), .ZN(n2262) );
  INVX0 U1417 ( .INP(n2295), .ZN(n2261) );
  INVX0 U1418 ( .INP(n2295), .ZN(n2260) );
  INVX0 U1419 ( .INP(n2295), .ZN(n2259) );
  INVX0 U1420 ( .INP(n2295), .ZN(n2258) );
  INVX0 U1421 ( .INP(n2296), .ZN(n2257) );
  INVX0 U1422 ( .INP(n2296), .ZN(n2256) );
  INVX0 U1423 ( .INP(n2296), .ZN(n2255) );
  INVX0 U1424 ( .INP(n2296), .ZN(n2254) );
  INVX0 U1425 ( .INP(n2296), .ZN(n2253) );
  INVX0 U1426 ( .INP(n2296), .ZN(n2252) );
  INVX0 U1427 ( .INP(n2296), .ZN(n2251) );
  INVX0 U1428 ( .INP(n2296), .ZN(n2250) );
  INVX0 U1429 ( .INP(n2296), .ZN(n2249) );
  INVX0 U1430 ( .INP(n2296), .ZN(n2248) );
  INVX0 U1431 ( .INP(n2296), .ZN(n2247) );
  INVX0 U1432 ( .INP(n2296), .ZN(n2246) );
  INVX0 U1433 ( .INP(n2297), .ZN(n2245) );
  INVX0 U1434 ( .INP(n2297), .ZN(n2244) );
  INVX0 U1435 ( .INP(n2297), .ZN(n2243) );
  INVX0 U1436 ( .INP(n2297), .ZN(n2242) );
  INVX0 U1437 ( .INP(n2297), .ZN(n2241) );
  INVX0 U1438 ( .INP(n2297), .ZN(n2240) );
  INVX0 U1439 ( .INP(n2297), .ZN(n2239) );
  INVX0 U1440 ( .INP(n2297), .ZN(n2238) );
  INVX0 U1441 ( .INP(n2297), .ZN(n2237) );
  INVX0 U1442 ( .INP(n2297), .ZN(n2236) );
  INVX0 U1443 ( .INP(n2297), .ZN(n2235) );
  INVX0 U1444 ( .INP(n2297), .ZN(n2234) );
  INVX0 U1445 ( .INP(n2298), .ZN(n2233) );
  INVX0 U1446 ( .INP(n2298), .ZN(n2232) );
  INVX0 U1447 ( .INP(n2298), .ZN(n2231) );
  INVX0 U1448 ( .INP(n2298), .ZN(n2230) );
  INVX0 U1449 ( .INP(n2298), .ZN(n2229) );
  INVX0 U1450 ( .INP(n2298), .ZN(n2228) );
  INVX0 U1451 ( .INP(n2298), .ZN(n2227) );
  INVX0 U1452 ( .INP(n2298), .ZN(n2226) );
  INVX0 U1453 ( .INP(n2298), .ZN(n2225) );
  INVX0 U1454 ( .INP(n2298), .ZN(n2224) );
  INVX0 U1455 ( .INP(n2298), .ZN(n2223) );
  INVX0 U1456 ( .INP(n2298), .ZN(n2222) );
  NAND2X1 U1457 ( .IN1(n2050), .IN2(\r[2][0] ), .QN(n2008) );
  NAND2X1 U1458 ( .IN1(n2050), .IN2(\r[2][1] ), .QN(n2004) );
  NAND2X1 U1459 ( .IN1(n2050), .IN2(\r[2][2] ), .QN(n2000) );
  NAND2X1 U1460 ( .IN1(n2050), .IN2(\r[2][3] ), .QN(n1996) );
  NAND2X1 U1461 ( .IN1(n2050), .IN2(\r[2][4] ), .QN(n1992) );
  NAND2X1 U1462 ( .IN1(n2050), .IN2(\r[2][5] ), .QN(n1988) );
  NAND2X1 U1463 ( .IN1(n2050), .IN2(\r[2][6] ), .QN(n1984) );
  NAND2X1 U1464 ( .IN1(n2050), .IN2(\r[2][7] ), .QN(n1980) );
  NAND2X1 U1465 ( .IN1(n2050), .IN2(\r[2][8] ), .QN(n1976) );
  NAND2X1 U1466 ( .IN1(n2050), .IN2(\r[2][9] ), .QN(n1972) );
  NAND2X1 U1467 ( .IN1(n2049), .IN2(\r[2][10] ), .QN(n1968) );
  NAND2X1 U1468 ( .IN1(n2050), .IN2(\r[2][11] ), .QN(n1964) );
  NAND2X1 U1469 ( .IN1(n2050), .IN2(\r[2][12] ), .QN(n1960) );
  NAND2X1 U1470 ( .IN1(n2050), .IN2(\r[2][13] ), .QN(n1956) );
  NAND2X1 U1471 ( .IN1(n2050), .IN2(\r[2][14] ), .QN(n1952) );
  NAND2X1 U1472 ( .IN1(n2050), .IN2(\r[2][15] ), .QN(n1948) );
  NAND2X1 U1473 ( .IN1(n2050), .IN2(\r[2][16] ), .QN(n1944) );
  NAND2X1 U1474 ( .IN1(n2050), .IN2(\r[2][17] ), .QN(n1940) );
  NAND2X1 U1475 ( .IN1(n2050), .IN2(\r[2][18] ), .QN(n1936) );
  NAND2X1 U1476 ( .IN1(n2049), .IN2(\r[2][19] ), .QN(n1932) );
  NAND2X1 U1477 ( .IN1(n2049), .IN2(\r[2][20] ), .QN(n1928) );
  NAND2X1 U1478 ( .IN1(n2050), .IN2(\r[2][21] ), .QN(n1924) );
  NAND2X1 U1479 ( .IN1(n2049), .IN2(\r[2][22] ), .QN(n1920) );
  NAND2X1 U1480 ( .IN1(n2049), .IN2(\r[2][23] ), .QN(n1916) );
  NAND2X1 U1481 ( .IN1(N17), .IN2(\r[2][24] ), .QN(n1912) );
  NAND2X1 U1482 ( .IN1(n2049), .IN2(\r[2][25] ), .QN(n1908) );
  NAND2X1 U1483 ( .IN1(n2049), .IN2(\r[2][26] ), .QN(n1904) );
  NAND2X1 U1484 ( .IN1(N17), .IN2(\r[2][27] ), .QN(n1900) );
  NAND2X1 U1485 ( .IN1(n2049), .IN2(\r[2][28] ), .QN(n1896) );
  NAND2X1 U1486 ( .IN1(n2049), .IN2(\r[2][29] ), .QN(n1892) );
  NAND2X1 U1487 ( .IN1(N17), .IN2(\r[2][30] ), .QN(n1888) );
  NAND2X1 U1488 ( .IN1(n2049), .IN2(\r[2][31] ), .QN(n1884) );
  NAND2X1 U1489 ( .IN1(n1558), .IN2(\r[2][0] ), .QN(n1516) );
  NAND2X1 U1490 ( .IN1(n1558), .IN2(\r[2][1] ), .QN(n1512) );
  NAND2X1 U1491 ( .IN1(n1558), .IN2(\r[2][2] ), .QN(n1508) );
  NAND2X1 U1492 ( .IN1(n1558), .IN2(\r[2][3] ), .QN(n1504) );
  NAND2X1 U1493 ( .IN1(n1558), .IN2(\r[2][4] ), .QN(n1500) );
  NAND2X1 U1494 ( .IN1(n1558), .IN2(\r[2][5] ), .QN(n1496) );
  NAND2X1 U1495 ( .IN1(n1558), .IN2(\r[2][6] ), .QN(n1492) );
  NAND2X1 U1496 ( .IN1(n1558), .IN2(\r[2][7] ), .QN(n1488) );
  NAND2X1 U1497 ( .IN1(n1558), .IN2(\r[2][8] ), .QN(n1484) );
  NAND2X1 U1498 ( .IN1(n1558), .IN2(\r[2][9] ), .QN(n1480) );
  NAND2X1 U1499 ( .IN1(n1557), .IN2(\r[2][10] ), .QN(n1476) );
  NAND2X1 U1500 ( .IN1(n1558), .IN2(\r[2][11] ), .QN(n1472) );
  NAND2X1 U1501 ( .IN1(n1558), .IN2(\r[2][12] ), .QN(n1468) );
  NAND2X1 U1502 ( .IN1(n1558), .IN2(\r[2][13] ), .QN(n1464) );
  NAND2X1 U1503 ( .IN1(n1558), .IN2(\r[2][14] ), .QN(n1460) );
  NAND2X1 U1504 ( .IN1(n1558), .IN2(\r[2][15] ), .QN(n1456) );
  NAND2X1 U1505 ( .IN1(n1558), .IN2(\r[2][16] ), .QN(n1452) );
  NAND2X1 U1506 ( .IN1(n1558), .IN2(\r[2][17] ), .QN(n1448) );
  NAND2X1 U1507 ( .IN1(n1558), .IN2(\r[2][18] ), .QN(n1444) );
  NAND2X1 U1508 ( .IN1(n1557), .IN2(\r[2][19] ), .QN(n1440) );
  NAND2X1 U1509 ( .IN1(n1557), .IN2(\r[2][20] ), .QN(n1436) );
  NAND2X1 U1510 ( .IN1(n1558), .IN2(\r[2][21] ), .QN(n1432) );
  NAND2X1 U1511 ( .IN1(n1557), .IN2(\r[2][22] ), .QN(n1428) );
  NAND2X1 U1512 ( .IN1(n1557), .IN2(\r[2][23] ), .QN(n1424) );
  NAND2X1 U1513 ( .IN1(N12), .IN2(\r[2][24] ), .QN(n1420) );
  NAND2X1 U1514 ( .IN1(n1557), .IN2(\r[2][25] ), .QN(n1416) );
  NAND2X1 U1515 ( .IN1(n1557), .IN2(\r[2][26] ), .QN(n1412) );
  NAND2X1 U1516 ( .IN1(N12), .IN2(\r[2][27] ), .QN(n1408) );
  NAND2X1 U1517 ( .IN1(n1557), .IN2(\r[2][28] ), .QN(n1404) );
  NAND2X1 U1518 ( .IN1(n1557), .IN2(\r[2][29] ), .QN(n1400) );
  NAND2X1 U1519 ( .IN1(N12), .IN2(\r[2][30] ), .QN(n1396) );
  NAND2X1 U1520 ( .IN1(n1557), .IN2(\r[2][31] ), .QN(n1392) );
  NAND2X1 U1521 ( .IN1(n2011), .IN2(n2010), .QN(n1572) );
  NAND2X1 U1522 ( .IN1(\r[1][0] ), .IN2(n2035), .QN(n2009) );
  NAND2X1 U1523 ( .IN1(n2007), .IN2(n2006), .QN(n1582) );
  NAND2X1 U1524 ( .IN1(\r[1][1] ), .IN2(n2035), .QN(n2005) );
  NAND2X1 U1525 ( .IN1(n2003), .IN2(n2002), .QN(n1592) );
  NAND2X1 U1526 ( .IN1(\r[1][2] ), .IN2(n2035), .QN(n2001) );
  NAND2X1 U1527 ( .IN1(n1999), .IN2(n1998), .QN(n1602) );
  NAND2X1 U1528 ( .IN1(\r[1][3] ), .IN2(n2035), .QN(n1997) );
  NAND2X1 U1529 ( .IN1(n1995), .IN2(n1994), .QN(n1612) );
  NAND2X1 U1530 ( .IN1(\r[1][4] ), .IN2(n2035), .QN(n1993) );
  NAND2X1 U1531 ( .IN1(n1991), .IN2(n1990), .QN(n1622) );
  NAND2X1 U1532 ( .IN1(\r[1][5] ), .IN2(n2035), .QN(n1989) );
  NAND2X1 U1533 ( .IN1(n1987), .IN2(n1986), .QN(n1632) );
  NAND2X1 U1534 ( .IN1(\r[1][6] ), .IN2(n2035), .QN(n1985) );
  NAND2X1 U1535 ( .IN1(n1983), .IN2(n1982), .QN(n1642) );
  NAND2X1 U1536 ( .IN1(\r[1][7] ), .IN2(n2035), .QN(n1981) );
  NAND2X1 U1537 ( .IN1(n1979), .IN2(n1978), .QN(n1652) );
  NAND2X1 U1538 ( .IN1(\r[1][8] ), .IN2(n2036), .QN(n1977) );
  NAND2X1 U1539 ( .IN1(n1975), .IN2(n1974), .QN(n1662) );
  NAND2X1 U1540 ( .IN1(\r[1][9] ), .IN2(n2036), .QN(n1973) );
  NAND2X1 U1541 ( .IN1(n1971), .IN2(n1970), .QN(n1672) );
  NAND2X1 U1542 ( .IN1(\r[1][10] ), .IN2(n2036), .QN(n1969) );
  NAND2X1 U1543 ( .IN1(n1967), .IN2(n1966), .QN(n1682) );
  NAND2X1 U1544 ( .IN1(\r[1][11] ), .IN2(n2036), .QN(n1965) );
  NAND2X1 U1545 ( .IN1(n1963), .IN2(n1962), .QN(n1692) );
  NAND2X1 U1546 ( .IN1(\r[1][12] ), .IN2(n2036), .QN(n1961) );
  NAND2X1 U1547 ( .IN1(n1959), .IN2(n1958), .QN(n1702) );
  NAND2X1 U1548 ( .IN1(\r[1][13] ), .IN2(n2036), .QN(n1957) );
  NAND2X1 U1549 ( .IN1(n1955), .IN2(n1954), .QN(n1712) );
  NAND2X1 U1550 ( .IN1(\r[1][14] ), .IN2(n2036), .QN(n1953) );
  NAND2X1 U1551 ( .IN1(n1951), .IN2(n1950), .QN(n1722) );
  NAND2X1 U1552 ( .IN1(\r[1][15] ), .IN2(n2036), .QN(n1949) );
  NAND2X1 U1553 ( .IN1(n1947), .IN2(n1946), .QN(n1732) );
  NAND2X1 U1554 ( .IN1(\r[1][16] ), .IN2(n2036), .QN(n1945) );
  NAND2X1 U1555 ( .IN1(n1943), .IN2(n1942), .QN(n1742) );
  NAND2X1 U1556 ( .IN1(\r[1][17] ), .IN2(n2036), .QN(n1941) );
  NAND2X1 U1557 ( .IN1(n1939), .IN2(n1938), .QN(n1752) );
  NAND2X1 U1558 ( .IN1(\r[1][18] ), .IN2(n2036), .QN(n1937) );
  NAND2X1 U1559 ( .IN1(n1935), .IN2(n1934), .QN(n1762) );
  NAND2X1 U1560 ( .IN1(\r[1][19] ), .IN2(n2036), .QN(n1933) );
  NAND2X1 U1561 ( .IN1(n1931), .IN2(n1930), .QN(n1772) );
  NAND2X1 U1562 ( .IN1(\r[1][20] ), .IN2(n2037), .QN(n1929) );
  NAND2X1 U1563 ( .IN1(n1927), .IN2(n1926), .QN(n1782) );
  NAND2X1 U1564 ( .IN1(\r[1][21] ), .IN2(n2037), .QN(n1925) );
  NAND2X1 U1565 ( .IN1(n1923), .IN2(n1922), .QN(n1792) );
  NAND2X1 U1566 ( .IN1(\r[1][22] ), .IN2(n2037), .QN(n1921) );
  NAND2X1 U1567 ( .IN1(n1919), .IN2(n1918), .QN(n1802) );
  NAND2X1 U1568 ( .IN1(\r[1][23] ), .IN2(n2037), .QN(n1917) );
  NAND2X1 U1569 ( .IN1(n1915), .IN2(n1914), .QN(n1812) );
  NAND2X1 U1570 ( .IN1(\r[1][24] ), .IN2(n2037), .QN(n1913) );
  NAND2X1 U1571 ( .IN1(n1911), .IN2(n1910), .QN(n1822) );
  NAND2X1 U1572 ( .IN1(\r[1][25] ), .IN2(n2037), .QN(n1909) );
  NAND2X1 U1573 ( .IN1(n1907), .IN2(n1906), .QN(n1832) );
  NAND2X1 U1574 ( .IN1(\r[1][26] ), .IN2(n2037), .QN(n1905) );
  NAND2X1 U1575 ( .IN1(n1903), .IN2(n1902), .QN(n1842) );
  NAND2X1 U1576 ( .IN1(\r[1][27] ), .IN2(n2037), .QN(n1901) );
  NAND2X1 U1577 ( .IN1(n1899), .IN2(n1898), .QN(n1852) );
  NAND2X1 U1578 ( .IN1(\r[1][28] ), .IN2(n2037), .QN(n1897) );
  NAND2X1 U1579 ( .IN1(n1895), .IN2(n1894), .QN(n1862) );
  NAND2X1 U1580 ( .IN1(\r[1][29] ), .IN2(n2037), .QN(n1893) );
  NAND2X1 U1581 ( .IN1(n1891), .IN2(n1890), .QN(n1872) );
  NAND2X1 U1582 ( .IN1(\r[1][30] ), .IN2(n2037), .QN(n1889) );
  NAND2X1 U1583 ( .IN1(n1887), .IN2(n1886), .QN(n1882) );
  NAND2X1 U1584 ( .IN1(\r[1][31] ), .IN2(n2037), .QN(n1885) );
  NAND2X1 U1585 ( .IN1(n1519), .IN2(n1518), .QN(n1080) );
  NAND2X1 U1586 ( .IN1(\r[1][0] ), .IN2(n1543), .QN(n1517) );
  NAND2X1 U1587 ( .IN1(n1515), .IN2(n1514), .QN(n1090) );
  NAND2X1 U1588 ( .IN1(\r[1][1] ), .IN2(n1543), .QN(n1513) );
  NAND2X1 U1589 ( .IN1(n1511), .IN2(n1510), .QN(n1100) );
  NAND2X1 U1590 ( .IN1(\r[1][2] ), .IN2(n1543), .QN(n1509) );
  NAND2X1 U1591 ( .IN1(n1507), .IN2(n1506), .QN(n1110) );
  NAND2X1 U1592 ( .IN1(\r[1][3] ), .IN2(n1543), .QN(n1505) );
  NAND2X1 U1593 ( .IN1(n1503), .IN2(n1502), .QN(n1120) );
  NAND2X1 U1594 ( .IN1(\r[1][4] ), .IN2(n1543), .QN(n1501) );
  NAND2X1 U1595 ( .IN1(n1499), .IN2(n1498), .QN(n1130) );
  NAND2X1 U1596 ( .IN1(\r[1][5] ), .IN2(n1543), .QN(n1497) );
  NAND2X1 U1597 ( .IN1(n1495), .IN2(n1494), .QN(n1140) );
  NAND2X1 U1598 ( .IN1(\r[1][6] ), .IN2(n1543), .QN(n1493) );
  NAND2X1 U1599 ( .IN1(n1491), .IN2(n1490), .QN(n1150) );
  NAND2X1 U1600 ( .IN1(\r[1][7] ), .IN2(n1543), .QN(n1489) );
  NAND2X1 U1601 ( .IN1(n1487), .IN2(n1486), .QN(n1160) );
  NAND2X1 U1602 ( .IN1(\r[1][8] ), .IN2(n1544), .QN(n1485) );
  NAND2X1 U1603 ( .IN1(n1483), .IN2(n1482), .QN(n1170) );
  NAND2X1 U1604 ( .IN1(\r[1][9] ), .IN2(n1544), .QN(n1481) );
  NAND2X1 U1605 ( .IN1(n1479), .IN2(n1478), .QN(n1180) );
  NAND2X1 U1606 ( .IN1(\r[1][10] ), .IN2(n1544), .QN(n1477) );
  NAND2X1 U1607 ( .IN1(n1475), .IN2(n1474), .QN(n1190) );
  NAND2X1 U1608 ( .IN1(\r[1][11] ), .IN2(n1544), .QN(n1473) );
  NAND2X1 U1609 ( .IN1(n1471), .IN2(n1470), .QN(n1200) );
  NAND2X1 U1610 ( .IN1(\r[1][12] ), .IN2(n1544), .QN(n1469) );
  NAND2X1 U1611 ( .IN1(n1467), .IN2(n1466), .QN(n1210) );
  NAND2X1 U1612 ( .IN1(\r[1][13] ), .IN2(n1544), .QN(n1465) );
  NAND2X1 U1613 ( .IN1(n1463), .IN2(n1462), .QN(n1220) );
  NAND2X1 U1614 ( .IN1(\r[1][14] ), .IN2(n1544), .QN(n1461) );
  NAND2X1 U1615 ( .IN1(n1459), .IN2(n1458), .QN(n1230) );
  NAND2X1 U1616 ( .IN1(\r[1][15] ), .IN2(n1544), .QN(n1457) );
  NAND2X1 U1617 ( .IN1(n1455), .IN2(n1454), .QN(n1240) );
  NAND2X1 U1618 ( .IN1(\r[1][16] ), .IN2(n1544), .QN(n1453) );
  NAND2X1 U1619 ( .IN1(n1451), .IN2(n1450), .QN(n1250) );
  NAND2X1 U1620 ( .IN1(\r[1][17] ), .IN2(n1544), .QN(n1449) );
  NAND2X1 U1621 ( .IN1(n1447), .IN2(n1446), .QN(n1260) );
  NAND2X1 U1622 ( .IN1(\r[1][18] ), .IN2(n1544), .QN(n1445) );
  NAND2X1 U1623 ( .IN1(n1443), .IN2(n1442), .QN(n1270) );
  NAND2X1 U1624 ( .IN1(\r[1][19] ), .IN2(n1544), .QN(n1441) );
  NAND2X1 U1625 ( .IN1(n1439), .IN2(n1438), .QN(n1280) );
  NAND2X1 U1626 ( .IN1(\r[1][20] ), .IN2(n1545), .QN(n1437) );
  NAND2X1 U1627 ( .IN1(n1435), .IN2(n1434), .QN(n1290) );
  NAND2X1 U1628 ( .IN1(\r[1][21] ), .IN2(n1545), .QN(n1433) );
  NAND2X1 U1629 ( .IN1(n1431), .IN2(n1430), .QN(n1300) );
  NAND2X1 U1630 ( .IN1(\r[1][22] ), .IN2(n1545), .QN(n1429) );
  NAND2X1 U1631 ( .IN1(n1427), .IN2(n1426), .QN(n1310) );
  NAND2X1 U1632 ( .IN1(\r[1][23] ), .IN2(n1545), .QN(n1425) );
  NAND2X1 U1633 ( .IN1(n1423), .IN2(n1422), .QN(n1320) );
  NAND2X1 U1634 ( .IN1(\r[1][24] ), .IN2(n1545), .QN(n1421) );
  NAND2X1 U1635 ( .IN1(n1419), .IN2(n1418), .QN(n1330) );
  NAND2X1 U1636 ( .IN1(\r[1][25] ), .IN2(n1545), .QN(n1417) );
  NAND2X1 U1637 ( .IN1(n1415), .IN2(n1414), .QN(n1340) );
  NAND2X1 U1638 ( .IN1(\r[1][26] ), .IN2(n1545), .QN(n1413) );
  NAND2X1 U1639 ( .IN1(n1411), .IN2(n1410), .QN(n1350) );
  NAND2X1 U1640 ( .IN1(\r[1][27] ), .IN2(n1545), .QN(n1409) );
  NAND2X1 U1641 ( .IN1(n1407), .IN2(n1406), .QN(n1360) );
  NAND2X1 U1642 ( .IN1(\r[1][28] ), .IN2(n1545), .QN(n1405) );
  NAND2X1 U1643 ( .IN1(n1403), .IN2(n1402), .QN(n1370) );
  NAND2X1 U1644 ( .IN1(\r[1][29] ), .IN2(n1545), .QN(n1401) );
  NAND2X1 U1645 ( .IN1(n1399), .IN2(n1398), .QN(n1380) );
  NAND2X1 U1646 ( .IN1(\r[1][30] ), .IN2(n1545), .QN(n1397) );
  NAND2X1 U1647 ( .IN1(n1395), .IN2(n1394), .QN(n1390) );
  NAND2X1 U1648 ( .IN1(\r[1][31] ), .IN2(n1545), .QN(n1393) );
  INVX0 U1649 ( .INP(N17), .ZN(n2036) );
  INVX0 U1650 ( .INP(N17), .ZN(n2037) );
  INVX0 U1651 ( .INP(N12), .ZN(n1544) );
  INVX0 U1652 ( .INP(N12), .ZN(n1545) );
  INVX0 U1653 ( .INP(wr_addr[2]), .ZN(n2301) );
  INVX0 U1654 ( .INP(wr_addr[1]), .ZN(n2302) );
  INVX0 U1655 ( .INP(wr_addr[0]), .ZN(n2303) );
  INVX0 U1656 ( .INP(wr_addr[4]), .ZN(n2299) );
  INVX0 U1657 ( .INP(wr_addr[3]), .ZN(n2300) );
  INVX0 U1658 ( .INP(nrst), .ZN(n2293) );
  INVX0 U1659 ( .INP(nrst), .ZN(n2294) );
  INVX0 U1660 ( .INP(nrst), .ZN(n2295) );
  INVX0 U1661 ( .INP(nrst), .ZN(n2296) );
  INVX0 U1662 ( .INP(nrst), .ZN(n2297) );
  INVX0 U1663 ( .INP(nrst), .ZN(n2298) );
  MUX41X1 U1664 ( .IN1(\r[28][0] ), .IN3(\r[30][0] ), .IN2(\r[29][0] ), .IN4(
        \r[31][0] ), .S0(n1547), .S1(n1525), .Q(n1072) );
  MUX41X1 U1665 ( .IN1(\r[24][0] ), .IN3(\r[26][0] ), .IN2(\r[25][0] ), .IN4(
        \r[27][0] ), .S0(n1557), .S1(n1542), .Q(n1073) );
  MUX41X1 U1666 ( .IN1(\r[20][0] ), .IN3(\r[22][0] ), .IN2(\r[21][0] ), .IN4(
        \r[23][0] ), .S0(n1551), .S1(n1522), .Q(n1074) );
  MUX41X1 U1667 ( .IN1(\r[16][0] ), .IN3(\r[18][0] ), .IN2(\r[17][0] ), .IN4(
        \r[19][0] ), .S0(n1551), .S1(n1522), .Q(n1075) );
  MUX41X1 U1668 ( .IN1(n1075), .IN3(n1073), .IN2(n1074), .IN4(n1072), .S0(N14),
        .S1(n1563), .Q(n1076) );
  MUX41X1 U1669 ( .IN1(\r[12][0] ), .IN3(\r[14][0] ), .IN2(\r[13][0] ), .IN4(
        \r[15][0] ), .S0(n1551), .S1(N11), .Q(n1077) );
  MUX41X1 U1670 ( .IN1(\r[8][0] ), .IN3(\r[10][0] ), .IN2(\r[9][0] ), .IN4(
        \r[11][0] ), .S0(n1551), .S1(N11), .Q(n1078) );
  MUX41X1 U1671 ( .IN1(\r[4][0] ), .IN3(\r[6][0] ), .IN2(\r[5][0] ), .IN4(
        \r[7][0] ), .S0(n1551), .S1(N11), .Q(n1079) );
  MUX41X1 U1672 ( .IN1(n1080), .IN3(n1078), .IN2(n1079), .IN4(n1077), .S0(N14),
        .S1(n1563), .Q(n1081) );
  MUX21X1 U1673 ( .IN1(n1081), .IN2(n1076), .S(N15), .Q(rd_dataA[0]) );
  MUX41X1 U1674 ( .IN1(\r[28][1] ), .IN3(\r[30][1] ), .IN2(\r[29][1] ), .IN4(
        \r[31][1] ), .S0(n1551), .S1(N11), .Q(n1082) );
  MUX41X1 U1675 ( .IN1(\r[24][1] ), .IN3(\r[26][1] ), .IN2(\r[25][1] ), .IN4(
        \r[27][1] ), .S0(n1551), .S1(N11), .Q(n1083) );
  MUX41X1 U1676 ( .IN1(\r[20][1] ), .IN3(\r[22][1] ), .IN2(\r[21][1] ), .IN4(
        \r[23][1] ), .S0(n1551), .S1(N11), .Q(n1084) );
  MUX41X1 U1677 ( .IN1(\r[16][1] ), .IN3(\r[18][1] ), .IN2(\r[17][1] ), .IN4(
        \r[19][1] ), .S0(n1551), .S1(n1522), .Q(n1085) );
  MUX41X1 U1678 ( .IN1(n1085), .IN3(n1083), .IN2(n1084), .IN4(n1082), .S0(N14),
        .S1(n1563), .Q(n1086) );
  MUX41X1 U1679 ( .IN1(\r[12][1] ), .IN3(\r[14][1] ), .IN2(\r[13][1] ), .IN4(
        \r[15][1] ), .S0(n1552), .S1(N11), .Q(n1087) );
  MUX41X1 U1680 ( .IN1(\r[8][1] ), .IN3(\r[10][1] ), .IN2(\r[9][1] ), .IN4(
        \r[11][1] ), .S0(n1552), .S1(N11), .Q(n1088) );
  MUX41X1 U1681 ( .IN1(\r[4][1] ), .IN3(\r[6][1] ), .IN2(\r[5][1] ), .IN4(
        \r[7][1] ), .S0(n1552), .S1(n1532), .Q(n1089) );
  MUX41X1 U1682 ( .IN1(n1090), .IN3(n1088), .IN2(n1089), .IN4(n1087), .S0(N14),
        .S1(n1563), .Q(n1091) );
  MUX21X1 U1683 ( .IN1(n1091), .IN2(n1086), .S(N15), .Q(rd_dataA[1]) );
  MUX41X1 U1684 ( .IN1(\r[28][2] ), .IN3(\r[30][2] ), .IN2(\r[29][2] ), .IN4(
        \r[31][2] ), .S0(n1552), .S1(n1532), .Q(n1092) );
  MUX41X1 U1685 ( .IN1(\r[24][2] ), .IN3(\r[26][2] ), .IN2(\r[25][2] ), .IN4(
        \r[27][2] ), .S0(n1552), .S1(n1532), .Q(n1093) );
  MUX41X1 U1686 ( .IN1(\r[20][2] ), .IN3(\r[22][2] ), .IN2(\r[21][2] ), .IN4(
        \r[23][2] ), .S0(n1552), .S1(n1532), .Q(n1094) );
  MUX41X1 U1687 ( .IN1(\r[16][2] ), .IN3(\r[18][2] ), .IN2(\r[17][2] ), .IN4(
        \r[19][2] ), .S0(n1552), .S1(n1532), .Q(n1095) );
  MUX41X1 U1688 ( .IN1(n1095), .IN3(n1093), .IN2(n1094), .IN4(n1092), .S0(N14),
        .S1(n1563), .Q(n1096) );
  MUX41X1 U1689 ( .IN1(\r[12][2] ), .IN3(\r[14][2] ), .IN2(\r[13][2] ), .IN4(
        \r[15][2] ), .S0(n1552), .S1(n1532), .Q(n1097) );
  MUX41X1 U1690 ( .IN1(\r[8][2] ), .IN3(\r[10][2] ), .IN2(\r[9][2] ), .IN4(
        \r[11][2] ), .S0(n1552), .S1(n1532), .Q(n1098) );
  MUX41X1 U1691 ( .IN1(\r[4][2] ), .IN3(\r[6][2] ), .IN2(\r[5][2] ), .IN4(
        \r[7][2] ), .S0(n1552), .S1(n1532), .Q(n1099) );
  MUX41X1 U1692 ( .IN1(n1100), .IN3(n1098), .IN2(n1099), .IN4(n1097), .S0(N14),
        .S1(n1563), .Q(n1101) );
  MUX21X1 U1693 ( .IN1(n1101), .IN2(n1096), .S(N15), .Q(rd_dataA[2]) );
  MUX41X1 U1694 ( .IN1(\r[28][3] ), .IN3(\r[30][3] ), .IN2(\r[29][3] ), .IN4(
        \r[31][3] ), .S0(n1552), .S1(n1532), .Q(n1102) );
  MUX41X1 U1695 ( .IN1(\r[24][3] ), .IN3(\r[26][3] ), .IN2(\r[25][3] ), .IN4(
        \r[27][3] ), .S0(n1552), .S1(n1532), .Q(n1103) );
  MUX41X1 U1696 ( .IN1(\r[20][3] ), .IN3(\r[22][3] ), .IN2(\r[21][3] ), .IN4(
        \r[23][3] ), .S0(n1552), .S1(n1532), .Q(n1104) );
  MUX41X1 U1697 ( .IN1(\r[16][3] ), .IN3(\r[18][3] ), .IN2(\r[17][3] ), .IN4(
        \r[19][3] ), .S0(n1552), .S1(n1532), .Q(n1105) );
  MUX41X1 U1698 ( .IN1(n1105), .IN3(n1103), .IN2(n1104), .IN4(n1102), .S0(N14),
        .S1(n1563), .Q(n1106) );
  MUX41X1 U1699 ( .IN1(\r[12][3] ), .IN3(\r[14][3] ), .IN2(\r[13][3] ), .IN4(
        \r[15][3] ), .S0(n1552), .S1(n1533), .Q(n1107) );
  MUX41X1 U1700 ( .IN1(\r[8][3] ), .IN3(\r[10][3] ), .IN2(\r[9][3] ), .IN4(
        \r[11][3] ), .S0(n1552), .S1(n1533), .Q(n1108) );
  MUX41X1 U1701 ( .IN1(\r[4][3] ), .IN3(\r[6][3] ), .IN2(\r[5][3] ), .IN4(
        \r[7][3] ), .S0(n1552), .S1(n1533), .Q(n1109) );
  MUX41X1 U1702 ( .IN1(n1110), .IN3(n1108), .IN2(n1109), .IN4(n1107), .S0(N14),
        .S1(n1563), .Q(n1111) );
  MUX21X1 U1703 ( .IN1(n1111), .IN2(n1106), .S(N15), .Q(rd_dataA[3]) );
  MUX41X1 U1704 ( .IN1(\r[28][4] ), .IN3(\r[30][4] ), .IN2(\r[29][4] ), .IN4(
        \r[31][4] ), .S0(n1552), .S1(n1533), .Q(n1112) );
  MUX41X1 U1705 ( .IN1(\r[24][4] ), .IN3(\r[26][4] ), .IN2(\r[25][4] ), .IN4(
        \r[27][4] ), .S0(n1552), .S1(n1533), .Q(n1113) );
  MUX41X1 U1706 ( .IN1(\r[20][4] ), .IN3(\r[22][4] ), .IN2(\r[21][4] ), .IN4(
        \r[23][4] ), .S0(n1552), .S1(n1533), .Q(n1114) );
  MUX41X1 U1707 ( .IN1(\r[16][4] ), .IN3(\r[18][4] ), .IN2(\r[17][4] ), .IN4(
        \r[19][4] ), .S0(n1552), .S1(n1533), .Q(n1115) );
  MUX41X1 U1708 ( .IN1(n1115), .IN3(n1113), .IN2(n1114), .IN4(n1112), .S0(N14),
        .S1(n1563), .Q(n1116) );
  MUX41X1 U1709 ( .IN1(\r[12][4] ), .IN3(\r[14][4] ), .IN2(\r[13][4] ), .IN4(
        \r[15][4] ), .S0(n1552), .S1(n1533), .Q(n1117) );
  MUX41X1 U1710 ( .IN1(\r[8][4] ), .IN3(\r[10][4] ), .IN2(\r[9][4] ), .IN4(
        \r[11][4] ), .S0(n1553), .S1(n1533), .Q(n1118) );
  MUX41X1 U1711 ( .IN1(\r[4][4] ), .IN3(\r[6][4] ), .IN2(\r[5][4] ), .IN4(
        \r[7][4] ), .S0(n1553), .S1(n1533), .Q(n1119) );
  MUX41X1 U1712 ( .IN1(n1120), .IN3(n1118), .IN2(n1119), .IN4(n1117), .S0(N14),
        .S1(n1563), .Q(n1121) );
  MUX21X1 U1713 ( .IN1(n1121), .IN2(n1116), .S(N15), .Q(rd_dataA[4]) );
  MUX41X1 U1714 ( .IN1(\r[28][5] ), .IN3(\r[30][5] ), .IN2(\r[29][5] ), .IN4(
        \r[31][5] ), .S0(n1553), .S1(n1533), .Q(n1122) );
  MUX41X1 U1715 ( .IN1(\r[24][5] ), .IN3(\r[26][5] ), .IN2(\r[25][5] ), .IN4(
        \r[27][5] ), .S0(n1553), .S1(n1533), .Q(n1123) );
  MUX41X1 U1716 ( .IN1(\r[20][5] ), .IN3(\r[22][5] ), .IN2(\r[21][5] ), .IN4(
        \r[23][5] ), .S0(n1553), .S1(n1534), .Q(n1124) );
  MUX41X1 U1717 ( .IN1(\r[16][5] ), .IN3(\r[18][5] ), .IN2(\r[17][5] ), .IN4(
        \r[19][5] ), .S0(n1553), .S1(n1534), .Q(n1125) );
  MUX41X1 U1718 ( .IN1(n1125), .IN3(n1123), .IN2(n1124), .IN4(n1122), .S0(N14),
        .S1(n1563), .Q(n1126) );
  MUX41X1 U1719 ( .IN1(\r[12][5] ), .IN3(\r[14][5] ), .IN2(\r[13][5] ), .IN4(
        \r[15][5] ), .S0(n1553), .S1(n1534), .Q(n1127) );
  MUX41X1 U1720 ( .IN1(\r[8][5] ), .IN3(\r[10][5] ), .IN2(\r[9][5] ), .IN4(
        \r[11][5] ), .S0(n1553), .S1(n1534), .Q(n1128) );
  MUX41X1 U1721 ( .IN1(\r[4][5] ), .IN3(\r[6][5] ), .IN2(\r[5][5] ), .IN4(
        \r[7][5] ), .S0(n1553), .S1(n1534), .Q(n1129) );
  MUX41X1 U1722 ( .IN1(n1130), .IN3(n1128), .IN2(n1129), .IN4(n1127), .S0(N14),
        .S1(n1563), .Q(n1131) );
  MUX21X1 U1723 ( .IN1(n1131), .IN2(n1126), .S(N15), .Q(rd_dataA[5]) );
  MUX41X1 U1724 ( .IN1(\r[28][6] ), .IN3(\r[30][6] ), .IN2(\r[29][6] ), .IN4(
        \r[31][6] ), .S0(n1553), .S1(n1534), .Q(n1132) );
  MUX41X1 U1725 ( .IN1(\r[24][6] ), .IN3(\r[26][6] ), .IN2(\r[25][6] ), .IN4(
        \r[27][6] ), .S0(n1553), .S1(n1534), .Q(n1133) );
  MUX41X1 U1726 ( .IN1(\r[20][6] ), .IN3(\r[22][6] ), .IN2(\r[21][6] ), .IN4(
        \r[23][6] ), .S0(n1553), .S1(n1534), .Q(n1134) );
  MUX41X1 U1727 ( .IN1(\r[16][6] ), .IN3(\r[18][6] ), .IN2(\r[17][6] ), .IN4(
        \r[19][6] ), .S0(n1553), .S1(n1534), .Q(n1135) );
  MUX41X1 U1728 ( .IN1(n1135), .IN3(n1133), .IN2(n1134), .IN4(n1132), .S0(N14),
        .S1(n1562), .Q(n1136) );
  MUX41X1 U1729 ( .IN1(\r[12][6] ), .IN3(\r[14][6] ), .IN2(\r[13][6] ), .IN4(
        \r[15][6] ), .S0(n1553), .S1(n1534), .Q(n1137) );
  MUX41X1 U1730 ( .IN1(\r[8][6] ), .IN3(\r[10][6] ), .IN2(\r[9][6] ), .IN4(
        \r[11][6] ), .S0(n1553), .S1(n1534), .Q(n1138) );
  MUX41X1 U1731 ( .IN1(\r[4][6] ), .IN3(\r[6][6] ), .IN2(\r[5][6] ), .IN4(
        \r[7][6] ), .S0(n1553), .S1(n1534), .Q(n1139) );
  MUX41X1 U1732 ( .IN1(n1140), .IN3(n1138), .IN2(n1139), .IN4(n1137), .S0(N14),
        .S1(n1562), .Q(n1141) );
  MUX21X1 U1733 ( .IN1(n1141), .IN2(n1136), .S(N15), .Q(rd_dataA[6]) );
  MUX41X1 U1734 ( .IN1(\r[28][7] ), .IN3(\r[30][7] ), .IN2(\r[29][7] ), .IN4(
        \r[31][7] ), .S0(n1553), .S1(n1535), .Q(n1142) );
  MUX41X1 U1735 ( .IN1(\r[24][7] ), .IN3(\r[26][7] ), .IN2(\r[25][7] ), .IN4(
        \r[27][7] ), .S0(n1553), .S1(n1535), .Q(n1143) );
  MUX41X1 U1736 ( .IN1(\r[20][7] ), .IN3(\r[22][7] ), .IN2(\r[21][7] ), .IN4(
        \r[23][7] ), .S0(n1553), .S1(n1535), .Q(n1144) );
  MUX41X1 U1737 ( .IN1(\r[16][7] ), .IN3(\r[18][7] ), .IN2(\r[17][7] ), .IN4(
        \r[19][7] ), .S0(n1553), .S1(n1535), .Q(n1145) );
  MUX41X1 U1738 ( .IN1(n1145), .IN3(n1143), .IN2(n1144), .IN4(n1142), .S0(N14),
        .S1(n1562), .Q(n1146) );
  MUX41X1 U1739 ( .IN1(\r[12][7] ), .IN3(\r[14][7] ), .IN2(\r[13][7] ), .IN4(
        \r[15][7] ), .S0(n1553), .S1(n1535), .Q(n1147) );
  MUX41X1 U1740 ( .IN1(\r[8][7] ), .IN3(\r[10][7] ), .IN2(\r[9][7] ), .IN4(
        \r[11][7] ), .S0(n1553), .S1(n1535), .Q(n1148) );
  MUX41X1 U1741 ( .IN1(\r[4][7] ), .IN3(\r[6][7] ), .IN2(\r[5][7] ), .IN4(
        \r[7][7] ), .S0(n1554), .S1(n1535), .Q(n1149) );
  MUX41X1 U1742 ( .IN1(n1150), .IN3(n1148), .IN2(n1149), .IN4(n1147), .S0(N14),
        .S1(n1562), .Q(n1151) );
  MUX21X1 U1743 ( .IN1(n1151), .IN2(n1146), .S(N15), .Q(rd_dataA[7]) );
  MUX41X1 U1744 ( .IN1(\r[28][8] ), .IN3(\r[30][8] ), .IN2(\r[29][8] ), .IN4(
        \r[31][8] ), .S0(n1554), .S1(n1535), .Q(n1152) );
  MUX41X1 U1745 ( .IN1(\r[24][8] ), .IN3(\r[26][8] ), .IN2(\r[25][8] ), .IN4(
        \r[27][8] ), .S0(n1554), .S1(n1535), .Q(n1153) );
  MUX41X1 U1746 ( .IN1(\r[20][8] ), .IN3(\r[22][8] ), .IN2(\r[21][8] ), .IN4(
        \r[23][8] ), .S0(n1554), .S1(n1535), .Q(n1154) );
  MUX41X1 U1747 ( .IN1(\r[16][8] ), .IN3(\r[18][8] ), .IN2(\r[17][8] ), .IN4(
        \r[19][8] ), .S0(n1554), .S1(n1535), .Q(n1155) );
  MUX41X1 U1748 ( .IN1(n1155), .IN3(n1153), .IN2(n1154), .IN4(n1152), .S0(N14),
        .S1(n1562), .Q(n1156) );
  MUX41X1 U1749 ( .IN1(\r[12][8] ), .IN3(\r[14][8] ), .IN2(\r[13][8] ), .IN4(
        \r[15][8] ), .S0(n1554), .S1(n1535), .Q(n1157) );
  MUX41X1 U1750 ( .IN1(\r[8][8] ), .IN3(\r[10][8] ), .IN2(\r[9][8] ), .IN4(
        \r[11][8] ), .S0(n1554), .S1(n1536), .Q(n1158) );
  MUX41X1 U1751 ( .IN1(\r[4][8] ), .IN3(\r[6][8] ), .IN2(\r[5][8] ), .IN4(
        \r[7][8] ), .S0(n1554), .S1(n1536), .Q(n1159) );
  MUX41X1 U1752 ( .IN1(n1160), .IN3(n1158), .IN2(n1159), .IN4(n1157), .S0(N14),
        .S1(n1562), .Q(n1161) );
  MUX21X1 U1753 ( .IN1(n1161), .IN2(n1156), .S(N15), .Q(rd_dataA[8]) );
  MUX41X1 U1754 ( .IN1(\r[28][9] ), .IN3(\r[30][9] ), .IN2(\r[29][9] ), .IN4(
        \r[31][9] ), .S0(n1554), .S1(n1536), .Q(n1162) );
  MUX41X1 U1755 ( .IN1(\r[24][9] ), .IN3(\r[26][9] ), .IN2(\r[25][9] ), .IN4(
        \r[27][9] ), .S0(n1554), .S1(n1536), .Q(n1163) );
  MUX41X1 U1756 ( .IN1(\r[20][9] ), .IN3(\r[22][9] ), .IN2(\r[21][9] ), .IN4(
        \r[23][9] ), .S0(n1554), .S1(n1536), .Q(n1164) );
  MUX41X1 U1757 ( .IN1(\r[16][9] ), .IN3(\r[18][9] ), .IN2(\r[17][9] ), .IN4(
        \r[19][9] ), .S0(n1554), .S1(n1536), .Q(n1165) );
  MUX41X1 U1758 ( .IN1(n1165), .IN3(n1163), .IN2(n1164), .IN4(n1162), .S0(N14),
        .S1(n1562), .Q(n1166) );
  MUX41X1 U1759 ( .IN1(\r[12][9] ), .IN3(\r[14][9] ), .IN2(\r[13][9] ), .IN4(
        \r[15][9] ), .S0(n1554), .S1(n1536), .Q(n1167) );
  MUX41X1 U1760 ( .IN1(\r[8][9] ), .IN3(\r[10][9] ), .IN2(\r[9][9] ), .IN4(
        \r[11][9] ), .S0(n1554), .S1(n1536), .Q(n1168) );
  MUX41X1 U1761 ( .IN1(\r[4][9] ), .IN3(\r[6][9] ), .IN2(\r[5][9] ), .IN4(
        \r[7][9] ), .S0(n1554), .S1(n1536), .Q(n1169) );
  MUX41X1 U1762 ( .IN1(n1170), .IN3(n1168), .IN2(n1169), .IN4(n1167), .S0(N14),
        .S1(n1562), .Q(n1171) );
  MUX21X1 U1763 ( .IN1(n1171), .IN2(n1166), .S(N15), .Q(rd_dataA[9]) );
  MUX41X1 U1764 ( .IN1(\r[28][10] ), .IN3(\r[30][10] ), .IN2(\r[29][10] ),
        .IN4(\r[31][10] ), .S0(n1554), .S1(n1536), .Q(n1172) );
  MUX41X1 U1765 ( .IN1(\r[24][10] ), .IN3(\r[26][10] ), .IN2(\r[25][10] ),
        .IN4(\r[27][10] ), .S0(n1554), .S1(n1536), .Q(n1173) );
  MUX41X1 U1766 ( .IN1(\r[20][10] ), .IN3(\r[22][10] ), .IN2(\r[21][10] ),
        .IN4(\r[23][10] ), .S0(n1554), .S1(n1536), .Q(n1174) );
  MUX41X1 U1767 ( .IN1(\r[16][10] ), .IN3(\r[18][10] ), .IN2(\r[17][10] ),
        .IN4(\r[19][10] ), .S0(n1554), .S1(n1537), .Q(n1175) );
  MUX41X1 U1768 ( .IN1(n1175), .IN3(n1173), .IN2(n1174), .IN4(n1172), .S0(N14),
        .S1(n1562), .Q(n1176) );
  MUX41X1 U1769 ( .IN1(\r[12][10] ), .IN3(\r[14][10] ), .IN2(\r[13][10] ),
        .IN4(\r[15][10] ), .S0(n1554), .S1(n1537), .Q(n1177) );
  MUX41X1 U1770 ( .IN1(\r[8][10] ), .IN3(\r[10][10] ), .IN2(\r[9][10] ), .IN4(
        \r[11][10] ), .S0(n1554), .S1(n1537), .Q(n1178) );
  MUX41X1 U1771 ( .IN1(\r[4][10] ), .IN3(\r[6][10] ), .IN2(\r[5][10] ), .IN4(
        \r[7][10] ), .S0(n1555), .S1(n1537), .Q(n1179) );
  MUX41X1 U1772 ( .IN1(n1180), .IN3(n1178), .IN2(n1179), .IN4(n1177), .S0(N14),
        .S1(n1562), .Q(n1181) );
  MUX21X1 U1773 ( .IN1(n1181), .IN2(n1176), .S(N15), .Q(rd_dataA[10]) );
  MUX41X1 U1774 ( .IN1(\r[28][11] ), .IN3(\r[30][11] ), .IN2(\r[29][11] ),
        .IN4(\r[31][11] ), .S0(n1555), .S1(n1537), .Q(n1182) );
  MUX41X1 U1775 ( .IN1(\r[24][11] ), .IN3(\r[26][11] ), .IN2(\r[25][11] ),
        .IN4(\r[27][11] ), .S0(n1555), .S1(n1537), .Q(n1183) );
  MUX41X1 U1776 ( .IN1(\r[20][11] ), .IN3(\r[22][11] ), .IN2(\r[21][11] ),
        .IN4(\r[23][11] ), .S0(n1555), .S1(n1537), .Q(n1184) );
  MUX41X1 U1777 ( .IN1(\r[16][11] ), .IN3(\r[18][11] ), .IN2(\r[17][11] ),
        .IN4(\r[19][11] ), .S0(n1555), .S1(n1537), .Q(n1185) );
  MUX41X1 U1778 ( .IN1(n1185), .IN3(n1183), .IN2(n1184), .IN4(n1182), .S0(N14),
        .S1(n1562), .Q(n1186) );
  MUX41X1 U1779 ( .IN1(\r[12][11] ), .IN3(\r[14][11] ), .IN2(\r[13][11] ),
        .IN4(\r[15][11] ), .S0(n1555), .S1(n1537), .Q(n1187) );
  MUX41X1 U1780 ( .IN1(\r[8][11] ), .IN3(\r[10][11] ), .IN2(\r[9][11] ), .IN4(
        \r[11][11] ), .S0(n1555), .S1(n1537), .Q(n1188) );
  MUX41X1 U1781 ( .IN1(\r[4][11] ), .IN3(\r[6][11] ), .IN2(\r[5][11] ), .IN4(
        \r[7][11] ), .S0(n1555), .S1(n1537), .Q(n1189) );
  MUX41X1 U1782 ( .IN1(n1190), .IN3(n1188), .IN2(n1189), .IN4(n1187), .S0(N14),
        .S1(n1562), .Q(n1191) );
  MUX21X1 U1783 ( .IN1(n1191), .IN2(n1186), .S(N15), .Q(rd_dataA[11]) );
  MUX41X1 U1784 ( .IN1(\r[28][12] ), .IN3(\r[30][12] ), .IN2(\r[29][12] ),
        .IN4(\r[31][12] ), .S0(n1555), .S1(n1538), .Q(n1192) );
  MUX41X1 U1785 ( .IN1(\r[24][12] ), .IN3(\r[26][12] ), .IN2(\r[25][12] ),
        .IN4(\r[27][12] ), .S0(n1555), .S1(n1538), .Q(n1193) );
  MUX41X1 U1786 ( .IN1(\r[20][12] ), .IN3(\r[22][12] ), .IN2(\r[21][12] ),
        .IN4(\r[23][12] ), .S0(n1555), .S1(n1538), .Q(n1194) );
  MUX41X1 U1787 ( .IN1(\r[16][12] ), .IN3(\r[18][12] ), .IN2(\r[17][12] ),
        .IN4(\r[19][12] ), .S0(n1555), .S1(n1538), .Q(n1195) );
  MUX41X1 U1788 ( .IN1(n1195), .IN3(n1193), .IN2(n1194), .IN4(n1192), .S0(N14),
        .S1(n1561), .Q(n1196) );
  MUX41X1 U1789 ( .IN1(\r[12][12] ), .IN3(\r[14][12] ), .IN2(\r[13][12] ),
        .IN4(\r[15][12] ), .S0(n1555), .S1(n1538), .Q(n1197) );
  MUX41X1 U1790 ( .IN1(\r[8][12] ), .IN3(\r[10][12] ), .IN2(\r[9][12] ), .IN4(
        \r[11][12] ), .S0(n1555), .S1(n1538), .Q(n1198) );
  MUX41X1 U1791 ( .IN1(\r[4][12] ), .IN3(\r[6][12] ), .IN2(\r[5][12] ), .IN4(
        \r[7][12] ), .S0(n1555), .S1(n1538), .Q(n1199) );
  MUX41X1 U1792 ( .IN1(n1200), .IN3(n1198), .IN2(n1199), .IN4(n1197), .S0(N14),
        .S1(n1561), .Q(n1201) );
  MUX21X1 U1793 ( .IN1(n1201), .IN2(n1196), .S(N15), .Q(rd_dataA[12]) );
  MUX41X1 U1794 ( .IN1(\r[28][13] ), .IN3(\r[30][13] ), .IN2(\r[29][13] ),
        .IN4(\r[31][13] ), .S0(n1555), .S1(n1538), .Q(n1202) );
  MUX41X1 U1795 ( .IN1(\r[24][13] ), .IN3(\r[26][13] ), .IN2(\r[25][13] ),
        .IN4(\r[27][13] ), .S0(n1555), .S1(n1538), .Q(n1203) );
  MUX41X1 U1796 ( .IN1(\r[20][13] ), .IN3(\r[22][13] ), .IN2(\r[21][13] ),
        .IN4(\r[23][13] ), .S0(n1555), .S1(n1538), .Q(n1204) );
  MUX41X1 U1797 ( .IN1(\r[16][13] ), .IN3(\r[18][13] ), .IN2(\r[17][13] ),
        .IN4(\r[19][13] ), .S0(n1555), .S1(n1538), .Q(n1205) );
  MUX41X1 U1798 ( .IN1(n1205), .IN3(n1203), .IN2(n1204), .IN4(n1202), .S0(N14),
        .S1(n1561), .Q(n1206) );
  MUX41X1 U1799 ( .IN1(\r[12][13] ), .IN3(\r[14][13] ), .IN2(\r[13][13] ),
        .IN4(\r[15][13] ), .S0(n1555), .S1(n1538), .Q(n1207) );
  MUX41X1 U1800 ( .IN1(\r[8][13] ), .IN3(\r[10][13] ), .IN2(\r[9][13] ), .IN4(
        \r[11][13] ), .S0(n1555), .S1(n1539), .Q(n1208) );
  MUX41X1 U1801 ( .IN1(\r[4][13] ), .IN3(\r[6][13] ), .IN2(\r[5][13] ), .IN4(
        \r[7][13] ), .S0(n1556), .S1(n1539), .Q(n1209) );
  MUX41X1 U1802 ( .IN1(n1210), .IN3(n1208), .IN2(n1209), .IN4(n1207), .S0(N14),
        .S1(n1561), .Q(n1211) );
  MUX21X1 U1803 ( .IN1(n1211), .IN2(n1206), .S(N15), .Q(rd_dataA[13]) );
  MUX41X1 U1804 ( .IN1(\r[28][14] ), .IN3(\r[30][14] ), .IN2(\r[29][14] ),
        .IN4(\r[31][14] ), .S0(n1555), .S1(n1539), .Q(n1212) );
  MUX41X1 U1805 ( .IN1(\r[24][14] ), .IN3(\r[26][14] ), .IN2(\r[25][14] ),
        .IN4(\r[27][14] ), .S0(n1556), .S1(n1539), .Q(n1213) );
  MUX41X1 U1806 ( .IN1(\r[20][14] ), .IN3(\r[22][14] ), .IN2(\r[21][14] ),
        .IN4(\r[23][14] ), .S0(n1556), .S1(n1539), .Q(n1214) );
  MUX41X1 U1807 ( .IN1(\r[16][14] ), .IN3(\r[18][14] ), .IN2(\r[17][14] ),
        .IN4(\r[19][14] ), .S0(n1556), .S1(n1539), .Q(n1215) );
  MUX41X1 U1808 ( .IN1(n1215), .IN3(n1213), .IN2(n1214), .IN4(n1212), .S0(N14),
        .S1(n1561), .Q(n1216) );
  MUX41X1 U1809 ( .IN1(\r[12][14] ), .IN3(\r[14][14] ), .IN2(\r[13][14] ),
        .IN4(\r[15][14] ), .S0(n1556), .S1(n1539), .Q(n1217) );
  MUX41X1 U1810 ( .IN1(\r[8][14] ), .IN3(\r[10][14] ), .IN2(\r[9][14] ), .IN4(
        \r[11][14] ), .S0(n1556), .S1(n1539), .Q(n1218) );
  MUX41X1 U1811 ( .IN1(\r[4][14] ), .IN3(\r[6][14] ), .IN2(\r[5][14] ), .IN4(
        \r[7][14] ), .S0(n1556), .S1(n1539), .Q(n1219) );
  MUX41X1 U1812 ( .IN1(n1220), .IN3(n1218), .IN2(n1219), .IN4(n1217), .S0(N14),
        .S1(n1561), .Q(n1221) );
  MUX21X1 U1813 ( .IN1(n1221), .IN2(n1216), .S(N15), .Q(rd_dataA[14]) );
  MUX41X1 U1814 ( .IN1(\r[28][15] ), .IN3(\r[30][15] ), .IN2(\r[29][15] ),
        .IN4(\r[31][15] ), .S0(n1556), .S1(n1539), .Q(n1222) );
  MUX41X1 U1815 ( .IN1(\r[24][15] ), .IN3(\r[26][15] ), .IN2(\r[25][15] ),
        .IN4(\r[27][15] ), .S0(n1556), .S1(n1539), .Q(n1223) );
  MUX41X1 U1816 ( .IN1(\r[20][15] ), .IN3(\r[22][15] ), .IN2(\r[21][15] ),
        .IN4(\r[23][15] ), .S0(n1556), .S1(n1539), .Q(n1224) );
  MUX41X1 U1817 ( .IN1(\r[16][15] ), .IN3(\r[18][15] ), .IN2(\r[17][15] ),
        .IN4(\r[19][15] ), .S0(n1556), .S1(n1540), .Q(n1225) );
  MUX41X1 U1818 ( .IN1(n1225), .IN3(n1223), .IN2(n1224), .IN4(n1222), .S0(N14),
        .S1(n1561), .Q(n1226) );
  MUX41X1 U1819 ( .IN1(\r[12][15] ), .IN3(\r[14][15] ), .IN2(\r[13][15] ),
        .IN4(\r[15][15] ), .S0(n1556), .S1(n1540), .Q(n1227) );
  MUX41X1 U1820 ( .IN1(\r[8][15] ), .IN3(\r[10][15] ), .IN2(\r[9][15] ), .IN4(
        \r[11][15] ), .S0(n1556), .S1(n1540), .Q(n1228) );
  MUX41X1 U1821 ( .IN1(\r[4][15] ), .IN3(\r[6][15] ), .IN2(\r[5][15] ), .IN4(
        \r[7][15] ), .S0(n1556), .S1(n1540), .Q(n1229) );
  MUX41X1 U1822 ( .IN1(n1230), .IN3(n1228), .IN2(n1229), .IN4(n1227), .S0(N14),
        .S1(n1561), .Q(n1231) );
  MUX21X1 U1823 ( .IN1(n1231), .IN2(n1226), .S(N15), .Q(rd_dataA[15]) );
  MUX41X1 U1824 ( .IN1(\r[28][16] ), .IN3(\r[30][16] ), .IN2(\r[29][16] ),
        .IN4(\r[31][16] ), .S0(n1556), .S1(n1540), .Q(n1232) );
  MUX41X1 U1825 ( .IN1(\r[24][16] ), .IN3(\r[26][16] ), .IN2(\r[25][16] ),
        .IN4(\r[27][16] ), .S0(n1556), .S1(n1540), .Q(n1233) );
  MUX41X1 U1826 ( .IN1(\r[20][16] ), .IN3(\r[22][16] ), .IN2(\r[21][16] ),
        .IN4(\r[23][16] ), .S0(n1556), .S1(n1540), .Q(n1234) );
  MUX41X1 U1827 ( .IN1(\r[16][16] ), .IN3(\r[18][16] ), .IN2(\r[17][16] ),
        .IN4(\r[19][16] ), .S0(n1557), .S1(n1540), .Q(n1235) );
  MUX41X1 U1828 ( .IN1(n1235), .IN3(n1233), .IN2(n1234), .IN4(n1232), .S0(N14),
        .S1(n1561), .Q(n1236) );
  MUX41X1 U1829 ( .IN1(\r[12][16] ), .IN3(\r[14][16] ), .IN2(\r[13][16] ),
        .IN4(\r[15][16] ), .S0(n1556), .S1(n1540), .Q(n1237) );
  MUX41X1 U1830 ( .IN1(\r[8][16] ), .IN3(\r[10][16] ), .IN2(\r[9][16] ), .IN4(
        \r[11][16] ), .S0(n1557), .S1(n1540), .Q(n1238) );
  MUX41X1 U1831 ( .IN1(\r[4][16] ), .IN3(\r[6][16] ), .IN2(\r[5][16] ), .IN4(
        \r[7][16] ), .S0(n1556), .S1(n1540), .Q(n1239) );
  MUX41X1 U1832 ( .IN1(n1240), .IN3(n1238), .IN2(n1239), .IN4(n1237), .S0(N14),
        .S1(n1561), .Q(n1241) );
  MUX21X1 U1833 ( .IN1(n1241), .IN2(n1236), .S(N15), .Q(rd_dataA[16]) );
  MUX41X1 U1834 ( .IN1(\r[28][17] ), .IN3(\r[30][17] ), .IN2(\r[29][17] ),
        .IN4(\r[31][17] ), .S0(n1556), .S1(n1540), .Q(n1242) );
  MUX41X1 U1835 ( .IN1(\r[24][17] ), .IN3(\r[26][17] ), .IN2(\r[25][17] ),
        .IN4(\r[27][17] ), .S0(n1557), .S1(n1541), .Q(n1243) );
  MUX41X1 U1836 ( .IN1(\r[20][17] ), .IN3(\r[22][17] ), .IN2(\r[21][17] ),
        .IN4(\r[23][17] ), .S0(n1557), .S1(n1541), .Q(n1244) );
  MUX41X1 U1837 ( .IN1(\r[16][17] ), .IN3(\r[18][17] ), .IN2(\r[17][17] ),
        .IN4(\r[19][17] ), .S0(n1556), .S1(n1541), .Q(n1245) );
  MUX41X1 U1838 ( .IN1(n1245), .IN3(n1243), .IN2(n1244), .IN4(n1242), .S0(N14),
        .S1(n1561), .Q(n1246) );
  MUX41X1 U1839 ( .IN1(\r[12][17] ), .IN3(\r[14][17] ), .IN2(\r[13][17] ),
        .IN4(\r[15][17] ), .S0(n1557), .S1(n1541), .Q(n1247) );
  MUX41X1 U1840 ( .IN1(\r[8][17] ), .IN3(\r[10][17] ), .IN2(\r[9][17] ), .IN4(
        \r[11][17] ), .S0(n1557), .S1(n1541), .Q(n1248) );
  MUX41X1 U1841 ( .IN1(\r[4][17] ), .IN3(\r[6][17] ), .IN2(\r[5][17] ), .IN4(
        \r[7][17] ), .S0(n1556), .S1(n1541), .Q(n1249) );
  MUX41X1 U1842 ( .IN1(n1250), .IN3(n1248), .IN2(n1249), .IN4(n1247), .S0(N14),
        .S1(n1561), .Q(n1251) );
  MUX21X1 U1843 ( .IN1(n1251), .IN2(n1246), .S(N15), .Q(rd_dataA[17]) );
  MUX41X1 U1844 ( .IN1(\r[28][18] ), .IN3(\r[30][18] ), .IN2(\r[29][18] ),
        .IN4(\r[31][18] ), .S0(n1557), .S1(n1541), .Q(n1252) );
  MUX41X1 U1845 ( .IN1(\r[24][18] ), .IN3(\r[26][18] ), .IN2(\r[25][18] ),
        .IN4(\r[27][18] ), .S0(n1554), .S1(n1541), .Q(n1253) );
  MUX41X1 U1846 ( .IN1(\r[20][18] ), .IN3(\r[22][18] ), .IN2(\r[21][18] ),
        .IN4(\r[23][18] ), .S0(n1547), .S1(n1541), .Q(n1254) );
  MUX41X1 U1847 ( .IN1(\r[16][18] ), .IN3(\r[18][18] ), .IN2(\r[17][18] ),
        .IN4(\r[19][18] ), .S0(n1547), .S1(n1541), .Q(n1255) );
  MUX41X1 U1848 ( .IN1(n1255), .IN3(n1253), .IN2(n1254), .IN4(n1252), .S0(N14),
        .S1(n1560), .Q(n1256) );
  MUX41X1 U1849 ( .IN1(\r[12][18] ), .IN3(\r[14][18] ), .IN2(\r[13][18] ),
        .IN4(\r[15][18] ), .S0(n1547), .S1(n1541), .Q(n1257) );
  MUX41X1 U1850 ( .IN1(\r[8][18] ), .IN3(\r[10][18] ), .IN2(\r[9][18] ), .IN4(
        \r[11][18] ), .S0(n1547), .S1(n1541), .Q(n1258) );
  MUX41X1 U1851 ( .IN1(\r[4][18] ), .IN3(\r[6][18] ), .IN2(\r[5][18] ), .IN4(
        \r[7][18] ), .S0(n1547), .S1(n1542), .Q(n1259) );
  MUX41X1 U1852 ( .IN1(n1260), .IN3(n1258), .IN2(n1259), .IN4(n1257), .S0(N14),
        .S1(n1560), .Q(n1261) );
  MUX21X1 U1853 ( .IN1(n1261), .IN2(n1256), .S(N15), .Q(rd_dataA[18]) );
  MUX41X1 U1854 ( .IN1(\r[28][19] ), .IN3(\r[30][19] ), .IN2(\r[29][19] ),
        .IN4(\r[31][19] ), .S0(n1547), .S1(n1542), .Q(n1262) );
  MUX41X1 U1855 ( .IN1(\r[24][19] ), .IN3(\r[26][19] ), .IN2(\r[25][19] ),
        .IN4(\r[27][19] ), .S0(n1547), .S1(n1542), .Q(n1263) );
  MUX41X1 U1856 ( .IN1(\r[20][19] ), .IN3(\r[22][19] ), .IN2(\r[21][19] ),
        .IN4(\r[23][19] ), .S0(n1547), .S1(n1542), .Q(n1264) );
  MUX41X1 U1857 ( .IN1(\r[16][19] ), .IN3(\r[18][19] ), .IN2(\r[17][19] ),
        .IN4(\r[19][19] ), .S0(n1547), .S1(n1542), .Q(n1265) );
  MUX41X1 U1858 ( .IN1(n1265), .IN3(n1263), .IN2(n1264), .IN4(n1262), .S0(N14),
        .S1(n1560), .Q(n1266) );
  MUX41X1 U1859 ( .IN1(\r[12][19] ), .IN3(\r[14][19] ), .IN2(\r[13][19] ),
        .IN4(\r[15][19] ), .S0(n1547), .S1(n1542), .Q(n1267) );
  MUX41X1 U1860 ( .IN1(\r[8][19] ), .IN3(\r[10][19] ), .IN2(\r[9][19] ), .IN4(
        \r[11][19] ), .S0(n1547), .S1(n1542), .Q(n1268) );
  MUX41X1 U1861 ( .IN1(\r[4][19] ), .IN3(\r[6][19] ), .IN2(\r[5][19] ), .IN4(
        \r[7][19] ), .S0(n1547), .S1(n1542), .Q(n1269) );
  MUX41X1 U1862 ( .IN1(n1270), .IN3(n1268), .IN2(n1269), .IN4(n1267), .S0(N14),
        .S1(n1560), .Q(n1271) );
  MUX21X1 U1863 ( .IN1(n1271), .IN2(n1266), .S(N15), .Q(rd_dataA[19]) );
  MUX41X1 U1864 ( .IN1(\r[28][20] ), .IN3(\r[30][20] ), .IN2(\r[29][20] ),
        .IN4(\r[31][20] ), .S0(n1547), .S1(n1542), .Q(n1272) );
  MUX41X1 U1865 ( .IN1(\r[24][20] ), .IN3(\r[26][20] ), .IN2(\r[25][20] ),
        .IN4(\r[27][20] ), .S0(n1547), .S1(n1542), .Q(n1273) );
  MUX41X1 U1866 ( .IN1(\r[20][20] ), .IN3(\r[22][20] ), .IN2(\r[21][20] ),
        .IN4(\r[23][20] ), .S0(n1547), .S1(n1542), .Q(n1274) );
  MUX41X1 U1867 ( .IN1(\r[16][20] ), .IN3(\r[18][20] ), .IN2(\r[17][20] ),
        .IN4(\r[19][20] ), .S0(n1547), .S1(n1537), .Q(n1275) );
  MUX41X1 U1868 ( .IN1(n1275), .IN3(n1273), .IN2(n1274), .IN4(n1272), .S0(N14),
        .S1(n1560), .Q(n1276) );
  MUX41X1 U1869 ( .IN1(\r[12][20] ), .IN3(\r[14][20] ), .IN2(\r[13][20] ),
        .IN4(\r[15][20] ), .S0(n1549), .S1(n1528), .Q(n1277) );
  MUX41X1 U1870 ( .IN1(\r[8][20] ), .IN3(\r[10][20] ), .IN2(\r[9][20] ), .IN4(
        \r[11][20] ), .S0(n1547), .S1(n1525), .Q(n1278) );
  MUX41X1 U1871 ( .IN1(\r[4][20] ), .IN3(\r[6][20] ), .IN2(\r[5][20] ), .IN4(
        \r[7][20] ), .S0(n1548), .S1(n1525), .Q(n1279) );
  MUX41X1 U1872 ( .IN1(n1280), .IN3(n1278), .IN2(n1279), .IN4(n1277), .S0(N14),
        .S1(n1560), .Q(n1281) );
  MUX21X1 U1873 ( .IN1(n1281), .IN2(n1276), .S(N15), .Q(rd_dataA[20]) );
  MUX41X1 U1874 ( .IN1(\r[28][21] ), .IN3(\r[30][21] ), .IN2(\r[29][21] ),
        .IN4(\r[31][21] ), .S0(n1548), .S1(n1525), .Q(n1282) );
  MUX41X1 U1875 ( .IN1(\r[24][21] ), .IN3(\r[26][21] ), .IN2(\r[25][21] ),
        .IN4(\r[27][21] ), .S0(n1548), .S1(n1525), .Q(n1283) );
  MUX41X1 U1876 ( .IN1(\r[20][21] ), .IN3(\r[22][21] ), .IN2(\r[21][21] ),
        .IN4(\r[23][21] ), .S0(n1548), .S1(n1525), .Q(n1284) );
  MUX41X1 U1877 ( .IN1(\r[16][21] ), .IN3(\r[18][21] ), .IN2(\r[17][21] ),
        .IN4(\r[19][21] ), .S0(n1548), .S1(n1525), .Q(n1285) );
  MUX41X1 U1878 ( .IN1(n1285), .IN3(n1283), .IN2(n1284), .IN4(n1282), .S0(N14),
        .S1(n1560), .Q(n1286) );
  MUX41X1 U1879 ( .IN1(\r[12][21] ), .IN3(\r[14][21] ), .IN2(\r[13][21] ),
        .IN4(\r[15][21] ), .S0(n1548), .S1(n1525), .Q(n1287) );
  MUX41X1 U1880 ( .IN1(\r[8][21] ), .IN3(\r[10][21] ), .IN2(\r[9][21] ), .IN4(
        \r[11][21] ), .S0(n1548), .S1(n1526), .Q(n1288) );
  MUX41X1 U1881 ( .IN1(\r[4][21] ), .IN3(\r[6][21] ), .IN2(\r[5][21] ), .IN4(
        \r[7][21] ), .S0(n1548), .S1(n1526), .Q(n1289) );
  MUX41X1 U1882 ( .IN1(n1290), .IN3(n1288), .IN2(n1289), .IN4(n1287), .S0(N14),
        .S1(n1560), .Q(n1291) );
  MUX21X1 U1883 ( .IN1(n1291), .IN2(n1286), .S(N15), .Q(rd_dataA[21]) );
  MUX41X1 U1884 ( .IN1(\r[28][22] ), .IN3(\r[30][22] ), .IN2(\r[29][22] ),
        .IN4(\r[31][22] ), .S0(n1548), .S1(n1526), .Q(n1292) );
  MUX41X1 U1885 ( .IN1(\r[24][22] ), .IN3(\r[26][22] ), .IN2(\r[25][22] ),
        .IN4(\r[27][22] ), .S0(n1548), .S1(n1526), .Q(n1293) );
  MUX41X1 U1886 ( .IN1(\r[20][22] ), .IN3(\r[22][22] ), .IN2(\r[21][22] ),
        .IN4(\r[23][22] ), .S0(n1548), .S1(n1526), .Q(n1294) );
  MUX41X1 U1887 ( .IN1(\r[16][22] ), .IN3(\r[18][22] ), .IN2(\r[17][22] ),
        .IN4(\r[19][22] ), .S0(n1548), .S1(n1526), .Q(n1295) );
  MUX41X1 U1888 ( .IN1(n1295), .IN3(n1293), .IN2(n1294), .IN4(n1292), .S0(N14),
        .S1(n1560), .Q(n1296) );
  MUX41X1 U1889 ( .IN1(\r[12][22] ), .IN3(\r[14][22] ), .IN2(\r[13][22] ),
        .IN4(\r[15][22] ), .S0(n1548), .S1(n1526), .Q(n1297) );
  MUX41X1 U1890 ( .IN1(\r[8][22] ), .IN3(\r[10][22] ), .IN2(\r[9][22] ), .IN4(
        \r[11][22] ), .S0(n1548), .S1(n1526), .Q(n1298) );
  MUX41X1 U1891 ( .IN1(\r[4][22] ), .IN3(\r[6][22] ), .IN2(\r[5][22] ), .IN4(
        \r[7][22] ), .S0(n1548), .S1(n1526), .Q(n1299) );
  MUX41X1 U1892 ( .IN1(n1300), .IN3(n1298), .IN2(n1299), .IN4(n1297), .S0(N14),
        .S1(n1560), .Q(n1301) );
  MUX21X1 U1893 ( .IN1(n1301), .IN2(n1296), .S(N15), .Q(rd_dataA[22]) );
  MUX41X1 U1894 ( .IN1(\r[28][23] ), .IN3(\r[30][23] ), .IN2(\r[29][23] ),
        .IN4(\r[31][23] ), .S0(n1548), .S1(n1526), .Q(n1302) );
  MUX41X1 U1895 ( .IN1(\r[24][23] ), .IN3(\r[26][23] ), .IN2(\r[25][23] ),
        .IN4(\r[27][23] ), .S0(n1548), .S1(n1526), .Q(n1303) );
  MUX41X1 U1896 ( .IN1(\r[20][23] ), .IN3(\r[22][23] ), .IN2(\r[21][23] ),
        .IN4(\r[23][23] ), .S0(n1548), .S1(n1526), .Q(n1304) );
  MUX41X1 U1897 ( .IN1(\r[16][23] ), .IN3(\r[18][23] ), .IN2(\r[17][23] ),
        .IN4(\r[19][23] ), .S0(n1548), .S1(n1527), .Q(n1305) );
  MUX41X1 U1898 ( .IN1(n1305), .IN3(n1303), .IN2(n1304), .IN4(n1302), .S0(N14),
        .S1(n1560), .Q(n1306) );
  MUX41X1 U1899 ( .IN1(\r[12][23] ), .IN3(\r[14][23] ), .IN2(\r[13][23] ),
        .IN4(\r[15][23] ), .S0(n1548), .S1(n1527), .Q(n1307) );
  MUX41X1 U1900 ( .IN1(\r[8][23] ), .IN3(\r[10][23] ), .IN2(\r[9][23] ), .IN4(
        \r[11][23] ), .S0(n1548), .S1(n1527), .Q(n1308) );
  MUX41X1 U1901 ( .IN1(\r[4][23] ), .IN3(\r[6][23] ), .IN2(\r[5][23] ), .IN4(
        \r[7][23] ), .S0(n1548), .S1(n1527), .Q(n1309) );
  MUX41X1 U1902 ( .IN1(n1310), .IN3(n1308), .IN2(n1309), .IN4(n1307), .S0(N14),
        .S1(n1560), .Q(n1311) );
  MUX21X1 U1903 ( .IN1(n1311), .IN2(n1306), .S(N15), .Q(rd_dataA[23]) );
  MUX41X1 U1904 ( .IN1(\r[28][24] ), .IN3(\r[30][24] ), .IN2(\r[29][24] ),
        .IN4(\r[31][24] ), .S0(n1549), .S1(n1527), .Q(n1312) );
  MUX41X1 U1905 ( .IN1(\r[24][24] ), .IN3(\r[26][24] ), .IN2(\r[25][24] ),
        .IN4(\r[27][24] ), .S0(n1549), .S1(n1527), .Q(n1313) );
  MUX41X1 U1906 ( .IN1(\r[20][24] ), .IN3(\r[22][24] ), .IN2(\r[21][24] ),
        .IN4(\r[23][24] ), .S0(n1549), .S1(n1527), .Q(n1314) );
  MUX41X1 U1907 ( .IN1(\r[16][24] ), .IN3(\r[18][24] ), .IN2(\r[17][24] ),
        .IN4(\r[19][24] ), .S0(n1549), .S1(n1527), .Q(n1315) );
  MUX41X1 U1908 ( .IN1(n1315), .IN3(n1313), .IN2(n1314), .IN4(n1312), .S0(N14),
        .S1(N13), .Q(n1316) );
  MUX41X1 U1909 ( .IN1(\r[12][24] ), .IN3(\r[14][24] ), .IN2(\r[13][24] ),
        .IN4(\r[15][24] ), .S0(n1549), .S1(n1527), .Q(n1317) );
  MUX41X1 U1910 ( .IN1(\r[8][24] ), .IN3(\r[10][24] ), .IN2(\r[9][24] ), .IN4(
        \r[11][24] ), .S0(n1549), .S1(n1527), .Q(n1318) );
  MUX41X1 U1911 ( .IN1(\r[4][24] ), .IN3(\r[6][24] ), .IN2(\r[5][24] ), .IN4(
        \r[7][24] ), .S0(n1549), .S1(n1527), .Q(n1319) );
  MUX41X1 U1912 ( .IN1(n1320), .IN3(n1318), .IN2(n1319), .IN4(n1317), .S0(N14),
        .S1(N13), .Q(n1321) );
  MUX21X1 U1913 ( .IN1(n1321), .IN2(n1316), .S(N15), .Q(rd_dataA[24]) );
  MUX41X1 U1914 ( .IN1(\r[28][25] ), .IN3(\r[30][25] ), .IN2(\r[29][25] ),
        .IN4(\r[31][25] ), .S0(n1549), .S1(n1527), .Q(n1322) );
  MUX41X1 U1915 ( .IN1(\r[24][25] ), .IN3(\r[26][25] ), .IN2(\r[25][25] ),
        .IN4(\r[27][25] ), .S0(n1549), .S1(n1528), .Q(n1323) );
  MUX41X1 U1916 ( .IN1(\r[20][25] ), .IN3(\r[22][25] ), .IN2(\r[21][25] ),
        .IN4(\r[23][25] ), .S0(n1549), .S1(n1528), .Q(n1324) );
  MUX41X1 U1917 ( .IN1(\r[16][25] ), .IN3(\r[18][25] ), .IN2(\r[17][25] ),
        .IN4(\r[19][25] ), .S0(n1549), .S1(n1528), .Q(n1325) );
  MUX41X1 U1918 ( .IN1(n1325), .IN3(n1323), .IN2(n1324), .IN4(n1322), .S0(N14),
        .S1(N13), .Q(n1326) );
  MUX41X1 U1919 ( .IN1(\r[12][25] ), .IN3(\r[14][25] ), .IN2(\r[13][25] ),
        .IN4(\r[15][25] ), .S0(n1549), .S1(n1528), .Q(n1327) );
  MUX41X1 U1920 ( .IN1(\r[8][25] ), .IN3(\r[10][25] ), .IN2(\r[9][25] ), .IN4(
        \r[11][25] ), .S0(n1549), .S1(n1528), .Q(n1328) );
  MUX41X1 U1921 ( .IN1(\r[4][25] ), .IN3(\r[6][25] ), .IN2(\r[5][25] ), .IN4(
        \r[7][25] ), .S0(n1549), .S1(n1528), .Q(n1329) );
  MUX41X1 U1922 ( .IN1(n1330), .IN3(n1328), .IN2(n1329), .IN4(n1327), .S0(N14),
        .S1(N13), .Q(n1331) );
  MUX21X1 U1923 ( .IN1(n1331), .IN2(n1326), .S(N15), .Q(rd_dataA[25]) );
  MUX41X1 U1924 ( .IN1(\r[28][26] ), .IN3(\r[30][26] ), .IN2(\r[29][26] ),
        .IN4(\r[31][26] ), .S0(n1549), .S1(n1528), .Q(n1332) );
  MUX41X1 U1925 ( .IN1(\r[24][26] ), .IN3(\r[26][26] ), .IN2(\r[25][26] ),
        .IN4(\r[27][26] ), .S0(n1549), .S1(n1528), .Q(n1333) );
  MUX41X1 U1926 ( .IN1(\r[20][26] ), .IN3(\r[22][26] ), .IN2(\r[21][26] ),
        .IN4(\r[23][26] ), .S0(n1549), .S1(n1528), .Q(n1334) );
  MUX41X1 U1927 ( .IN1(\r[16][26] ), .IN3(\r[18][26] ), .IN2(\r[17][26] ),
        .IN4(\r[19][26] ), .S0(n1549), .S1(n1528), .Q(n1335) );
  MUX41X1 U1928 ( .IN1(n1335), .IN3(n1333), .IN2(n1334), .IN4(n1332), .S0(N14),
        .S1(N13), .Q(n1336) );
  MUX41X1 U1929 ( .IN1(\r[12][26] ), .IN3(\r[14][26] ), .IN2(\r[13][26] ),
        .IN4(\r[15][26] ), .S0(n1549), .S1(n1528), .Q(n1337) );
  MUX41X1 U1930 ( .IN1(\r[8][26] ), .IN3(\r[10][26] ), .IN2(\r[9][26] ), .IN4(
        \r[11][26] ), .S0(n1549), .S1(n1529), .Q(n1338) );
  MUX41X1 U1931 ( .IN1(\r[4][26] ), .IN3(\r[6][26] ), .IN2(\r[5][26] ), .IN4(
        \r[7][26] ), .S0(n1549), .S1(n1529), .Q(n1339) );
  MUX41X1 U1932 ( .IN1(n1340), .IN3(n1338), .IN2(n1339), .IN4(n1337), .S0(N14),
        .S1(N13), .Q(n1341) );
  MUX21X1 U1933 ( .IN1(n1341), .IN2(n1336), .S(N15), .Q(rd_dataA[26]) );
  MUX41X1 U1934 ( .IN1(\r[28][27] ), .IN3(\r[30][27] ), .IN2(\r[29][27] ),
        .IN4(\r[31][27] ), .S0(n1550), .S1(n1529), .Q(n1342) );
  MUX41X1 U1935 ( .IN1(\r[24][27] ), .IN3(\r[26][27] ), .IN2(\r[25][27] ),
        .IN4(\r[27][27] ), .S0(n1550), .S1(n1529), .Q(n1343) );
  MUX41X1 U1936 ( .IN1(\r[20][27] ), .IN3(\r[22][27] ), .IN2(\r[21][27] ),
        .IN4(\r[23][27] ), .S0(n1550), .S1(n1529), .Q(n1344) );
  MUX41X1 U1937 ( .IN1(\r[16][27] ), .IN3(\r[18][27] ), .IN2(\r[17][27] ),
        .IN4(\r[19][27] ), .S0(n1550), .S1(n1529), .Q(n1345) );
  MUX41X1 U1938 ( .IN1(n1345), .IN3(n1343), .IN2(n1344), .IN4(n1342), .S0(N14),
        .S1(N13), .Q(n1346) );
  MUX41X1 U1939 ( .IN1(\r[12][27] ), .IN3(\r[14][27] ), .IN2(\r[13][27] ),
        .IN4(\r[15][27] ), .S0(n1550), .S1(n1529), .Q(n1347) );
  MUX41X1 U1940 ( .IN1(\r[8][27] ), .IN3(\r[10][27] ), .IN2(\r[9][27] ), .IN4(
        \r[11][27] ), .S0(n1550), .S1(n1529), .Q(n1348) );
  MUX41X1 U1941 ( .IN1(\r[4][27] ), .IN3(\r[6][27] ), .IN2(\r[5][27] ), .IN4(
        \r[7][27] ), .S0(n1550), .S1(n1529), .Q(n1349) );
  MUX41X1 U1942 ( .IN1(n1350), .IN3(n1348), .IN2(n1349), .IN4(n1347), .S0(N14),
        .S1(N13), .Q(n1351) );
  MUX21X1 U1943 ( .IN1(n1351), .IN2(n1346), .S(N15), .Q(rd_dataA[27]) );
  MUX41X1 U1944 ( .IN1(\r[28][28] ), .IN3(\r[30][28] ), .IN2(\r[29][28] ),
        .IN4(\r[31][28] ), .S0(n1550), .S1(n1529), .Q(n1352) );
  MUX41X1 U1945 ( .IN1(\r[24][28] ), .IN3(\r[26][28] ), .IN2(\r[25][28] ),
        .IN4(\r[27][28] ), .S0(n1550), .S1(n1529), .Q(n1353) );
  MUX41X1 U1946 ( .IN1(\r[20][28] ), .IN3(\r[22][28] ), .IN2(\r[21][28] ),
        .IN4(\r[23][28] ), .S0(n1550), .S1(n1529), .Q(n1354) );
  MUX41X1 U1947 ( .IN1(\r[16][28] ), .IN3(\r[18][28] ), .IN2(\r[17][28] ),
        .IN4(\r[19][28] ), .S0(n1550), .S1(n1530), .Q(n1355) );
  MUX41X1 U1948 ( .IN1(n1355), .IN3(n1353), .IN2(n1354), .IN4(n1352), .S0(N14),
        .S1(N13), .Q(n1356) );
  MUX41X1 U1949 ( .IN1(\r[12][28] ), .IN3(\r[14][28] ), .IN2(\r[13][28] ),
        .IN4(\r[15][28] ), .S0(n1550), .S1(n1530), .Q(n1357) );
  MUX41X1 U1950 ( .IN1(\r[8][28] ), .IN3(\r[10][28] ), .IN2(\r[9][28] ), .IN4(
        \r[11][28] ), .S0(n1550), .S1(n1530), .Q(n1358) );
  MUX41X1 U1951 ( .IN1(\r[4][28] ), .IN3(\r[6][28] ), .IN2(\r[5][28] ), .IN4(
        \r[7][28] ), .S0(n1550), .S1(n1530), .Q(n1359) );
  MUX41X1 U1952 ( .IN1(n1360), .IN3(n1358), .IN2(n1359), .IN4(n1357), .S0(N14),
        .S1(N13), .Q(n1361) );
  MUX21X1 U1953 ( .IN1(n1361), .IN2(n1356), .S(N15), .Q(rd_dataA[28]) );
  MUX41X1 U1954 ( .IN1(\r[28][29] ), .IN3(\r[30][29] ), .IN2(\r[29][29] ),
        .IN4(\r[31][29] ), .S0(n1550), .S1(n1530), .Q(n1362) );
  MUX41X1 U1955 ( .IN1(\r[24][29] ), .IN3(\r[26][29] ), .IN2(\r[25][29] ),
        .IN4(\r[27][29] ), .S0(n1550), .S1(n1530), .Q(n1363) );
  MUX41X1 U1956 ( .IN1(\r[20][29] ), .IN3(\r[22][29] ), .IN2(\r[21][29] ),
        .IN4(\r[23][29] ), .S0(n1550), .S1(n1530), .Q(n1364) );
  MUX41X1 U1957 ( .IN1(\r[16][29] ), .IN3(\r[18][29] ), .IN2(\r[17][29] ),
        .IN4(\r[19][29] ), .S0(n1550), .S1(n1530), .Q(n1365) );
  MUX41X1 U1958 ( .IN1(n1365), .IN3(n1363), .IN2(n1364), .IN4(n1362), .S0(N14),
        .S1(N13), .Q(n1366) );
  MUX41X1 U1959 ( .IN1(\r[12][29] ), .IN3(\r[14][29] ), .IN2(\r[13][29] ),
        .IN4(\r[15][29] ), .S0(n1550), .S1(n1530), .Q(n1367) );
  MUX41X1 U1960 ( .IN1(\r[8][29] ), .IN3(\r[10][29] ), .IN2(\r[9][29] ), .IN4(
        \r[11][29] ), .S0(n1550), .S1(n1530), .Q(n1368) );
  MUX41X1 U1961 ( .IN1(\r[4][29] ), .IN3(\r[6][29] ), .IN2(\r[5][29] ), .IN4(
        \r[7][29] ), .S0(n1550), .S1(n1530), .Q(n1369) );
  MUX41X1 U1962 ( .IN1(n1370), .IN3(n1368), .IN2(n1369), .IN4(n1367), .S0(N14),
        .S1(N13), .Q(n1371) );
  MUX21X1 U1963 ( .IN1(n1371), .IN2(n1366), .S(N15), .Q(rd_dataA[29]) );
  MUX41X1 U1964 ( .IN1(\r[28][30] ), .IN3(\r[30][30] ), .IN2(\r[29][30] ),
        .IN4(\r[31][30] ), .S0(n1550), .S1(n1530), .Q(n1372) );
  MUX41X1 U1965 ( .IN1(\r[24][30] ), .IN3(\r[26][30] ), .IN2(\r[25][30] ),
        .IN4(\r[27][30] ), .S0(n1551), .S1(n1531), .Q(n1373) );
  MUX41X1 U1966 ( .IN1(\r[20][30] ), .IN3(\r[22][30] ), .IN2(\r[21][30] ),
        .IN4(\r[23][30] ), .S0(n1551), .S1(n1531), .Q(n1374) );
  MUX41X1 U1967 ( .IN1(\r[16][30] ), .IN3(\r[18][30] ), .IN2(\r[17][30] ),
        .IN4(\r[19][30] ), .S0(n1551), .S1(n1531), .Q(n1375) );
  MUX41X1 U1968 ( .IN1(n1375), .IN3(n1373), .IN2(n1374), .IN4(n1372), .S0(N14),
        .S1(N13), .Q(n1376) );
  MUX41X1 U1969 ( .IN1(\r[12][30] ), .IN3(\r[14][30] ), .IN2(\r[13][30] ),
        .IN4(\r[15][30] ), .S0(n1551), .S1(n1531), .Q(n1377) );
  MUX41X1 U1970 ( .IN1(\r[8][30] ), .IN3(\r[10][30] ), .IN2(\r[9][30] ), .IN4(
        \r[11][30] ), .S0(n1551), .S1(n1531), .Q(n1378) );
  MUX41X1 U1971 ( .IN1(\r[4][30] ), .IN3(\r[6][30] ), .IN2(\r[5][30] ), .IN4(
        \r[7][30] ), .S0(n1551), .S1(n1531), .Q(n1379) );
  MUX41X1 U1972 ( .IN1(n1380), .IN3(n1378), .IN2(n1379), .IN4(n1377), .S0(N14),
        .S1(N13), .Q(n1381) );
  MUX21X1 U1973 ( .IN1(n1381), .IN2(n1376), .S(N15), .Q(rd_dataA[30]) );
  MUX41X1 U1974 ( .IN1(\r[28][31] ), .IN3(\r[30][31] ), .IN2(\r[29][31] ),
        .IN4(\r[31][31] ), .S0(n1551), .S1(n1531), .Q(n1382) );
  MUX41X1 U1975 ( .IN1(\r[24][31] ), .IN3(\r[26][31] ), .IN2(\r[25][31] ),
        .IN4(\r[27][31] ), .S0(n1551), .S1(n1531), .Q(n1383) );
  MUX41X1 U1976 ( .IN1(\r[20][31] ), .IN3(\r[22][31] ), .IN2(\r[21][31] ),
        .IN4(\r[23][31] ), .S0(n1551), .S1(n1531), .Q(n1384) );
  MUX41X1 U1977 ( .IN1(\r[16][31] ), .IN3(\r[18][31] ), .IN2(\r[17][31] ),
        .IN4(\r[19][31] ), .S0(n1551), .S1(n1531), .Q(n1385) );
  MUX41X1 U1978 ( .IN1(n1385), .IN3(n1383), .IN2(n1384), .IN4(n1382), .S0(N14),
        .S1(N13), .Q(n1386) );
  MUX41X1 U1979 ( .IN1(\r[12][31] ), .IN3(\r[14][31] ), .IN2(\r[13][31] ),
        .IN4(\r[15][31] ), .S0(n1551), .S1(n1531), .Q(n1387) );
  MUX41X1 U1980 ( .IN1(\r[8][31] ), .IN3(\r[10][31] ), .IN2(\r[9][31] ), .IN4(
        \r[11][31] ), .S0(n1551), .S1(n1531), .Q(n1388) );
  MUX41X1 U1981 ( .IN1(\r[4][31] ), .IN3(\r[6][31] ), .IN2(\r[5][31] ), .IN4(
        \r[7][31] ), .S0(n1551), .S1(N11), .Q(n1389) );
  MUX41X1 U1982 ( .IN1(n1390), .IN3(n1388), .IN2(n1389), .IN4(n1387), .S0(N14),
        .S1(N13), .Q(n1391) );
  MUX21X1 U1983 ( .IN1(n1391), .IN2(n1386), .S(N15), .Q(rd_dataA[31]) );
  MUX21X1 U1984 ( .IN1(n1392), .IN2(n1393), .S(n1525), .Q(n1395) );
  NAND3X0 U1985 ( .IN1(\r[3][31] ), .IN2(n1522), .IN3(n1547), .QN(n1394) );
  MUX21X1 U1986 ( .IN1(n1396), .IN2(n1397), .S(n1523), .Q(n1399) );
  NAND3X0 U1987 ( .IN1(\r[3][30] ), .IN2(n1522), .IN3(n1547), .QN(n1398) );
  MUX21X1 U1988 ( .IN1(n1400), .IN2(n1401), .S(n1523), .Q(n1403) );
  NAND3X0 U1989 ( .IN1(\r[3][29] ), .IN2(n1522), .IN3(n1547), .QN(n1402) );
  MUX21X1 U1990 ( .IN1(n1404), .IN2(n1405), .S(n1523), .Q(n1407) );
  NAND3X0 U1991 ( .IN1(\r[3][28] ), .IN2(n1522), .IN3(n1547), .QN(n1406) );
  MUX21X1 U1992 ( .IN1(n1408), .IN2(n1409), .S(n1523), .Q(n1411) );
  NAND3X0 U1993 ( .IN1(\r[3][27] ), .IN2(n1522), .IN3(n1546), .QN(n1410) );
  MUX21X1 U1994 ( .IN1(n1412), .IN2(n1413), .S(n1523), .Q(n1415) );
  NAND3X0 U1995 ( .IN1(\r[3][26] ), .IN2(n1522), .IN3(n1546), .QN(n1414) );
  MUX21X1 U1996 ( .IN1(n1416), .IN2(n1417), .S(n1523), .Q(n1419) );
  NAND3X0 U1997 ( .IN1(\r[3][25] ), .IN2(n1523), .IN3(n1546), .QN(n1418) );
  MUX21X1 U1998 ( .IN1(n1420), .IN2(n1421), .S(n1523), .Q(n1423) );
  NAND3X0 U1999 ( .IN1(\r[3][24] ), .IN2(n1522), .IN3(n1546), .QN(n1422) );
  MUX21X1 U2000 ( .IN1(n1424), .IN2(n1425), .S(n1523), .Q(n1427) );
  NAND3X0 U2001 ( .IN1(\r[3][23] ), .IN2(n1523), .IN3(n1546), .QN(n1426) );
  MUX21X1 U2002 ( .IN1(n1428), .IN2(n1429), .S(n1524), .Q(n1431) );
  NAND3X0 U2003 ( .IN1(\r[3][22] ), .IN2(n1523), .IN3(n1546), .QN(n1430) );
  MUX21X1 U2004 ( .IN1(n1432), .IN2(n1433), .S(n1524), .Q(n1435) );
  NAND3X0 U2005 ( .IN1(\r[3][21] ), .IN2(n1523), .IN3(n1546), .QN(n1434) );
  MUX21X1 U2006 ( .IN1(n1436), .IN2(n1437), .S(n1524), .Q(n1439) );
  NAND3X0 U2007 ( .IN1(\r[3][20] ), .IN2(n1523), .IN3(n1546), .QN(n1438) );
  MUX21X1 U2008 ( .IN1(n1440), .IN2(n1441), .S(n1524), .Q(n1443) );
  NAND3X0 U2009 ( .IN1(\r[3][19] ), .IN2(n1523), .IN3(n1546), .QN(n1442) );
  MUX21X1 U2010 ( .IN1(n1444), .IN2(n1445), .S(n1524), .Q(n1447) );
  NAND3X0 U2011 ( .IN1(\r[3][18] ), .IN2(n1523), .IN3(n1546), .QN(n1446) );
  MUX21X1 U2012 ( .IN1(n1448), .IN2(n1449), .S(n1524), .Q(n1451) );
  NAND3X0 U2013 ( .IN1(\r[3][17] ), .IN2(n1523), .IN3(n1546), .QN(n1450) );
  MUX21X1 U2014 ( .IN1(n1452), .IN2(n1453), .S(n1524), .Q(n1455) );
  NAND3X0 U2015 ( .IN1(\r[3][16] ), .IN2(n1523), .IN3(n1546), .QN(n1454) );
  MUX21X1 U2016 ( .IN1(n1456), .IN2(n1457), .S(n1524), .Q(n1459) );
  NAND3X0 U2017 ( .IN1(\r[3][15] ), .IN2(n1523), .IN3(n1546), .QN(n1458) );
  MUX21X1 U2018 ( .IN1(n1460), .IN2(n1461), .S(n1524), .Q(n1463) );
  NAND3X0 U2019 ( .IN1(\r[3][14] ), .IN2(n1523), .IN3(n1546), .QN(n1462) );
  MUX21X1 U2020 ( .IN1(n1464), .IN2(n1465), .S(n1524), .Q(n1467) );
  NAND3X0 U2021 ( .IN1(\r[3][13] ), .IN2(n1523), .IN3(n1546), .QN(n1466) );
  MUX21X1 U2022 ( .IN1(n1468), .IN2(n1469), .S(n1524), .Q(n1471) );
  NAND3X0 U2023 ( .IN1(\r[3][12] ), .IN2(n1522), .IN3(n1546), .QN(n1470) );
  MUX21X1 U2024 ( .IN1(n1472), .IN2(n1473), .S(n1524), .Q(n1475) );
  NAND3X0 U2025 ( .IN1(\r[3][11] ), .IN2(n1523), .IN3(n1546), .QN(n1474) );
  MUX21X1 U2026 ( .IN1(n1476), .IN2(n1477), .S(n1524), .Q(n1479) );
  NAND3X0 U2027 ( .IN1(\r[3][10] ), .IN2(n1522), .IN3(n1546), .QN(n1478) );
  MUX21X1 U2028 ( .IN1(n1480), .IN2(n1481), .S(n1524), .Q(n1483) );
  NAND3X0 U2029 ( .IN1(\r[3][9] ), .IN2(n1522), .IN3(n1546), .QN(n1482) );
  MUX21X1 U2030 ( .IN1(n1484), .IN2(n1485), .S(n1524), .Q(n1487) );
  NAND3X0 U2031 ( .IN1(\r[3][8] ), .IN2(n1522), .IN3(n1546), .QN(n1486) );
  MUX21X1 U2032 ( .IN1(n1488), .IN2(n1489), .S(n1524), .Q(n1491) );
  NAND3X0 U2033 ( .IN1(\r[3][7] ), .IN2(n1522), .IN3(n1546), .QN(n1490) );
  MUX21X1 U2034 ( .IN1(n1492), .IN2(n1493), .S(n1524), .Q(n1495) );
  NAND3X0 U2035 ( .IN1(\r[3][6] ), .IN2(n1522), .IN3(n1546), .QN(n1494) );
  MUX21X1 U2036 ( .IN1(n1496), .IN2(n1497), .S(n1524), .Q(n1499) );
  NAND3X0 U2037 ( .IN1(\r[3][5] ), .IN2(n1522), .IN3(n1546), .QN(n1498) );
  MUX21X1 U2038 ( .IN1(n1500), .IN2(n1501), .S(n1525), .Q(n1503) );
  NAND3X0 U2039 ( .IN1(\r[3][4] ), .IN2(n1522), .IN3(n1546), .QN(n1502) );
  MUX21X1 U2040 ( .IN1(n1504), .IN2(n1505), .S(n1525), .Q(n1507) );
  NAND3X0 U2041 ( .IN1(\r[3][3] ), .IN2(n1522), .IN3(n1546), .QN(n1506) );
  MUX21X1 U2042 ( .IN1(n1508), .IN2(n1509), .S(n1525), .Q(n1511) );
  NAND3X0 U2043 ( .IN1(\r[3][2] ), .IN2(n1522), .IN3(n1546), .QN(n1510) );
  MUX21X1 U2044 ( .IN1(n1512), .IN2(n1513), .S(n1525), .Q(n1515) );
  NAND3X0 U2045 ( .IN1(\r[3][1] ), .IN2(n1522), .IN3(n1546), .QN(n1514) );
  MUX21X1 U2046 ( .IN1(n1516), .IN2(n1517), .S(n1525), .Q(n1519) );
  NAND3X0 U2047 ( .IN1(\r[3][0] ), .IN2(n1523), .IN3(n1547), .QN(n1518) );
  MUX41X1 U2048 ( .IN1(\r[28][0] ), .IN3(\r[30][0] ), .IN2(\r[29][0] ), .IN4(
        \r[31][0] ), .S0(n2039), .S1(n2017), .Q(n1564) );
  MUX41X1 U2049 ( .IN1(\r[24][0] ), .IN3(\r[26][0] ), .IN2(\r[25][0] ), .IN4(
        \r[27][0] ), .S0(n2049), .S1(n2034), .Q(n1565) );
  MUX41X1 U2050 ( .IN1(\r[20][0] ), .IN3(\r[22][0] ), .IN2(\r[21][0] ), .IN4(
        \r[23][0] ), .S0(n2043), .S1(n2014), .Q(n1566) );
  MUX41X1 U2051 ( .IN1(\r[16][0] ), .IN3(\r[18][0] ), .IN2(\r[17][0] ), .IN4(
        \r[19][0] ), .S0(n2043), .S1(n2014), .Q(n1567) );
  MUX41X1 U2052 ( .IN1(n1567), .IN3(n1565), .IN2(n1566), .IN4(n1564), .S0(N19),
        .S1(n2055), .Q(n1568) );
  MUX41X1 U2053 ( .IN1(\r[12][0] ), .IN3(\r[14][0] ), .IN2(\r[13][0] ), .IN4(
        \r[15][0] ), .S0(n2043), .S1(N16), .Q(n1569) );
  MUX41X1 U2054 ( .IN1(\r[8][0] ), .IN3(\r[10][0] ), .IN2(\r[9][0] ), .IN4(
        \r[11][0] ), .S0(n2043), .S1(N16), .Q(n1570) );
  MUX41X1 U2055 ( .IN1(\r[4][0] ), .IN3(\r[6][0] ), .IN2(\r[5][0] ), .IN4(
        \r[7][0] ), .S0(n2043), .S1(N16), .Q(n1571) );
  MUX41X1 U2056 ( .IN1(n1572), .IN3(n1570), .IN2(n1571), .IN4(n1569), .S0(N19),
        .S1(n2055), .Q(n1573) );
  MUX21X1 U2057 ( .IN1(n1573), .IN2(n1568), .S(N20), .Q(rd_dataB[0]) );
  MUX41X1 U2058 ( .IN1(\r[28][1] ), .IN3(\r[30][1] ), .IN2(\r[29][1] ), .IN4(
        \r[31][1] ), .S0(n2043), .S1(N16), .Q(n1574) );
  MUX41X1 U2059 ( .IN1(\r[24][1] ), .IN3(\r[26][1] ), .IN2(\r[25][1] ), .IN4(
        \r[27][1] ), .S0(n2043), .S1(N16), .Q(n1575) );
  MUX41X1 U2060 ( .IN1(\r[20][1] ), .IN3(\r[22][1] ), .IN2(\r[21][1] ), .IN4(
        \r[23][1] ), .S0(n2043), .S1(N16), .Q(n1576) );
  MUX41X1 U2061 ( .IN1(\r[16][1] ), .IN3(\r[18][1] ), .IN2(\r[17][1] ), .IN4(
        \r[19][1] ), .S0(n2043), .S1(n2014), .Q(n1577) );
  MUX41X1 U2062 ( .IN1(n1577), .IN3(n1575), .IN2(n1576), .IN4(n1574), .S0(N19),
        .S1(n2055), .Q(n1578) );
  MUX41X1 U2063 ( .IN1(\r[12][1] ), .IN3(\r[14][1] ), .IN2(\r[13][1] ), .IN4(
        \r[15][1] ), .S0(n2044), .S1(N16), .Q(n1579) );
  MUX41X1 U2064 ( .IN1(\r[8][1] ), .IN3(\r[10][1] ), .IN2(\r[9][1] ), .IN4(
        \r[11][1] ), .S0(n2044), .S1(N16), .Q(n1580) );
  MUX41X1 U2065 ( .IN1(\r[4][1] ), .IN3(\r[6][1] ), .IN2(\r[5][1] ), .IN4(
        \r[7][1] ), .S0(n2044), .S1(n2024), .Q(n1581) );
  MUX41X1 U2066 ( .IN1(n1582), .IN3(n1580), .IN2(n1581), .IN4(n1579), .S0(N19),
        .S1(n2055), .Q(n1583) );
  MUX21X1 U2067 ( .IN1(n1583), .IN2(n1578), .S(N20), .Q(rd_dataB[1]) );
  MUX41X1 U2068 ( .IN1(\r[28][2] ), .IN3(\r[30][2] ), .IN2(\r[29][2] ), .IN4(
        \r[31][2] ), .S0(n2044), .S1(n2024), .Q(n1584) );
  MUX41X1 U2069 ( .IN1(\r[24][2] ), .IN3(\r[26][2] ), .IN2(\r[25][2] ), .IN4(
        \r[27][2] ), .S0(n2044), .S1(n2024), .Q(n1585) );
  MUX41X1 U2070 ( .IN1(\r[20][2] ), .IN3(\r[22][2] ), .IN2(\r[21][2] ), .IN4(
        \r[23][2] ), .S0(n2044), .S1(n2024), .Q(n1586) );
  MUX41X1 U2071 ( .IN1(\r[16][2] ), .IN3(\r[18][2] ), .IN2(\r[17][2] ), .IN4(
        \r[19][2] ), .S0(n2044), .S1(n2024), .Q(n1587) );
  MUX41X1 U2072 ( .IN1(n1587), .IN3(n1585), .IN2(n1586), .IN4(n1584), .S0(N19),
        .S1(n2055), .Q(n1588) );
  MUX41X1 U2073 ( .IN1(\r[12][2] ), .IN3(\r[14][2] ), .IN2(\r[13][2] ), .IN4(
        \r[15][2] ), .S0(n2044), .S1(n2024), .Q(n1589) );
  MUX41X1 U2074 ( .IN1(\r[8][2] ), .IN3(\r[10][2] ), .IN2(\r[9][2] ), .IN4(
        \r[11][2] ), .S0(n2044), .S1(n2024), .Q(n1590) );
  MUX41X1 U2075 ( .IN1(\r[4][2] ), .IN3(\r[6][2] ), .IN2(\r[5][2] ), .IN4(
        \r[7][2] ), .S0(n2044), .S1(n2024), .Q(n1591) );
  MUX41X1 U2076 ( .IN1(n1592), .IN3(n1590), .IN2(n1591), .IN4(n1589), .S0(N19),
        .S1(n2055), .Q(n1593) );
  MUX21X1 U2077 ( .IN1(n1593), .IN2(n1588), .S(N20), .Q(rd_dataB[2]) );
  MUX41X1 U2078 ( .IN1(\r[28][3] ), .IN3(\r[30][3] ), .IN2(\r[29][3] ), .IN4(
        \r[31][3] ), .S0(n2044), .S1(n2024), .Q(n1594) );
  MUX41X1 U2079 ( .IN1(\r[24][3] ), .IN3(\r[26][3] ), .IN2(\r[25][3] ), .IN4(
        \r[27][3] ), .S0(n2044), .S1(n2024), .Q(n1595) );
  MUX41X1 U2080 ( .IN1(\r[20][3] ), .IN3(\r[22][3] ), .IN2(\r[21][3] ), .IN4(
        \r[23][3] ), .S0(n2044), .S1(n2024), .Q(n1596) );
  MUX41X1 U2081 ( .IN1(\r[16][3] ), .IN3(\r[18][3] ), .IN2(\r[17][3] ), .IN4(
        \r[19][3] ), .S0(n2044), .S1(n2024), .Q(n1597) );
  MUX41X1 U2082 ( .IN1(n1597), .IN3(n1595), .IN2(n1596), .IN4(n1594), .S0(N19),
        .S1(n2055), .Q(n1598) );
  MUX41X1 U2083 ( .IN1(\r[12][3] ), .IN3(\r[14][3] ), .IN2(\r[13][3] ), .IN4(
        \r[15][3] ), .S0(n2044), .S1(n2025), .Q(n1599) );
  MUX41X1 U2084 ( .IN1(\r[8][3] ), .IN3(\r[10][3] ), .IN2(\r[9][3] ), .IN4(
        \r[11][3] ), .S0(n2044), .S1(n2025), .Q(n1600) );
  MUX41X1 U2085 ( .IN1(\r[4][3] ), .IN3(\r[6][3] ), .IN2(\r[5][3] ), .IN4(
        \r[7][3] ), .S0(n2044), .S1(n2025), .Q(n1601) );
  MUX41X1 U2086 ( .IN1(n1602), .IN3(n1600), .IN2(n1601), .IN4(n1599), .S0(N19),
        .S1(n2055), .Q(n1603) );
  MUX21X1 U2087 ( .IN1(n1603), .IN2(n1598), .S(N20), .Q(rd_dataB[3]) );
  MUX41X1 U2088 ( .IN1(\r[28][4] ), .IN3(\r[30][4] ), .IN2(\r[29][4] ), .IN4(
        \r[31][4] ), .S0(n2044), .S1(n2025), .Q(n1604) );
  MUX41X1 U2089 ( .IN1(\r[24][4] ), .IN3(\r[26][4] ), .IN2(\r[25][4] ), .IN4(
        \r[27][4] ), .S0(n2044), .S1(n2025), .Q(n1605) );
  MUX41X1 U2090 ( .IN1(\r[20][4] ), .IN3(\r[22][4] ), .IN2(\r[21][4] ), .IN4(
        \r[23][4] ), .S0(n2044), .S1(n2025), .Q(n1606) );
  MUX41X1 U2091 ( .IN1(\r[16][4] ), .IN3(\r[18][4] ), .IN2(\r[17][4] ), .IN4(
        \r[19][4] ), .S0(n2044), .S1(n2025), .Q(n1607) );
  MUX41X1 U2092 ( .IN1(n1607), .IN3(n1605), .IN2(n1606), .IN4(n1604), .S0(N19),
        .S1(n2055), .Q(n1608) );
  MUX41X1 U2093 ( .IN1(\r[12][4] ), .IN3(\r[14][4] ), .IN2(\r[13][4] ), .IN4(
        \r[15][4] ), .S0(n2044), .S1(n2025), .Q(n1609) );
  MUX41X1 U2094 ( .IN1(\r[8][4] ), .IN3(\r[10][4] ), .IN2(\r[9][4] ), .IN4(
        \r[11][4] ), .S0(n2045), .S1(n2025), .Q(n1610) );
  MUX41X1 U2095 ( .IN1(\r[4][4] ), .IN3(\r[6][4] ), .IN2(\r[5][4] ), .IN4(
        \r[7][4] ), .S0(n2045), .S1(n2025), .Q(n1611) );
  MUX41X1 U2096 ( .IN1(n1612), .IN3(n1610), .IN2(n1611), .IN4(n1609), .S0(N19),
        .S1(n2055), .Q(n1613) );
  MUX21X1 U2097 ( .IN1(n1613), .IN2(n1608), .S(N20), .Q(rd_dataB[4]) );
  MUX41X1 U2098 ( .IN1(\r[28][5] ), .IN3(\r[30][5] ), .IN2(\r[29][5] ), .IN4(
        \r[31][5] ), .S0(n2045), .S1(n2025), .Q(n1614) );
  MUX41X1 U2099 ( .IN1(\r[24][5] ), .IN3(\r[26][5] ), .IN2(\r[25][5] ), .IN4(
        \r[27][5] ), .S0(n2045), .S1(n2025), .Q(n1615) );
  MUX41X1 U2100 ( .IN1(\r[20][5] ), .IN3(\r[22][5] ), .IN2(\r[21][5] ), .IN4(
        \r[23][5] ), .S0(n2045), .S1(n2026), .Q(n1616) );
  MUX41X1 U2101 ( .IN1(\r[16][5] ), .IN3(\r[18][5] ), .IN2(\r[17][5] ), .IN4(
        \r[19][5] ), .S0(n2045), .S1(n2026), .Q(n1617) );
  MUX41X1 U2102 ( .IN1(n1617), .IN3(n1615), .IN2(n1616), .IN4(n1614), .S0(N19),
        .S1(n2055), .Q(n1618) );
  MUX41X1 U2103 ( .IN1(\r[12][5] ), .IN3(\r[14][5] ), .IN2(\r[13][5] ), .IN4(
        \r[15][5] ), .S0(n2045), .S1(n2026), .Q(n1619) );
  MUX41X1 U2104 ( .IN1(\r[8][5] ), .IN3(\r[10][5] ), .IN2(\r[9][5] ), .IN4(
        \r[11][5] ), .S0(n2045), .S1(n2026), .Q(n1620) );
  MUX41X1 U2105 ( .IN1(\r[4][5] ), .IN3(\r[6][5] ), .IN2(\r[5][5] ), .IN4(
        \r[7][5] ), .S0(n2045), .S1(n2026), .Q(n1621) );
  MUX41X1 U2106 ( .IN1(n1622), .IN3(n1620), .IN2(n1621), .IN4(n1619), .S0(N19),
        .S1(n2055), .Q(n1623) );
  MUX21X1 U2107 ( .IN1(n1623), .IN2(n1618), .S(N20), .Q(rd_dataB[5]) );
  MUX41X1 U2108 ( .IN1(\r[28][6] ), .IN3(\r[30][6] ), .IN2(\r[29][6] ), .IN4(
        \r[31][6] ), .S0(n2045), .S1(n2026), .Q(n1624) );
  MUX41X1 U2109 ( .IN1(\r[24][6] ), .IN3(\r[26][6] ), .IN2(\r[25][6] ), .IN4(
        \r[27][6] ), .S0(n2045), .S1(n2026), .Q(n1625) );
  MUX41X1 U2110 ( .IN1(\r[20][6] ), .IN3(\r[22][6] ), .IN2(\r[21][6] ), .IN4(
        \r[23][6] ), .S0(n2045), .S1(n2026), .Q(n1626) );
  MUX41X1 U2111 ( .IN1(\r[16][6] ), .IN3(\r[18][6] ), .IN2(\r[17][6] ), .IN4(
        \r[19][6] ), .S0(n2045), .S1(n2026), .Q(n1627) );
  MUX41X1 U2112 ( .IN1(n1627), .IN3(n1625), .IN2(n1626), .IN4(n1624), .S0(N19),
        .S1(n2054), .Q(n1628) );
  MUX41X1 U2113 ( .IN1(\r[12][6] ), .IN3(\r[14][6] ), .IN2(\r[13][6] ), .IN4(
        \r[15][6] ), .S0(n2045), .S1(n2026), .Q(n1629) );
  MUX41X1 U2114 ( .IN1(\r[8][6] ), .IN3(\r[10][6] ), .IN2(\r[9][6] ), .IN4(
        \r[11][6] ), .S0(n2045), .S1(n2026), .Q(n1630) );
  MUX41X1 U2115 ( .IN1(\r[4][6] ), .IN3(\r[6][6] ), .IN2(\r[5][6] ), .IN4(
        \r[7][6] ), .S0(n2045), .S1(n2026), .Q(n1631) );
  MUX41X1 U2116 ( .IN1(n1632), .IN3(n1630), .IN2(n1631), .IN4(n1629), .S0(N19),
        .S1(n2054), .Q(n1633) );
  MUX21X1 U2117 ( .IN1(n1633), .IN2(n1628), .S(N20), .Q(rd_dataB[6]) );
  MUX41X1 U2118 ( .IN1(\r[28][7] ), .IN3(\r[30][7] ), .IN2(\r[29][7] ), .IN4(
        \r[31][7] ), .S0(n2045), .S1(n2027), .Q(n1634) );
  MUX41X1 U2119 ( .IN1(\r[24][7] ), .IN3(\r[26][7] ), .IN2(\r[25][7] ), .IN4(
        \r[27][7] ), .S0(n2045), .S1(n2027), .Q(n1635) );
  MUX41X1 U2120 ( .IN1(\r[20][7] ), .IN3(\r[22][7] ), .IN2(\r[21][7] ), .IN4(
        \r[23][7] ), .S0(n2045), .S1(n2027), .Q(n1636) );
  MUX41X1 U2121 ( .IN1(\r[16][7] ), .IN3(\r[18][7] ), .IN2(\r[17][7] ), .IN4(
        \r[19][7] ), .S0(n2045), .S1(n2027), .Q(n1637) );
  MUX41X1 U2122 ( .IN1(n1637), .IN3(n1635), .IN2(n1636), .IN4(n1634), .S0(N19),
        .S1(n2054), .Q(n1638) );
  MUX41X1 U2123 ( .IN1(\r[12][7] ), .IN3(\r[14][7] ), .IN2(\r[13][7] ), .IN4(
        \r[15][7] ), .S0(n2045), .S1(n2027), .Q(n1639) );
  MUX41X1 U2124 ( .IN1(\r[8][7] ), .IN3(\r[10][7] ), .IN2(\r[9][7] ), .IN4(
        \r[11][7] ), .S0(n2045), .S1(n2027), .Q(n1640) );
  MUX41X1 U2125 ( .IN1(\r[4][7] ), .IN3(\r[6][7] ), .IN2(\r[5][7] ), .IN4(
        \r[7][7] ), .S0(n2046), .S1(n2027), .Q(n1641) );
  MUX41X1 U2126 ( .IN1(n1642), .IN3(n1640), .IN2(n1641), .IN4(n1639), .S0(N19),
        .S1(n2054), .Q(n1643) );
  MUX21X1 U2127 ( .IN1(n1643), .IN2(n1638), .S(N20), .Q(rd_dataB[7]) );
  MUX41X1 U2128 ( .IN1(\r[28][8] ), .IN3(\r[30][8] ), .IN2(\r[29][8] ), .IN4(
        \r[31][8] ), .S0(n2046), .S1(n2027), .Q(n1644) );
  MUX41X1 U2129 ( .IN1(\r[24][8] ), .IN3(\r[26][8] ), .IN2(\r[25][8] ), .IN4(
        \r[27][8] ), .S0(n2046), .S1(n2027), .Q(n1645) );
  MUX41X1 U2130 ( .IN1(\r[20][8] ), .IN3(\r[22][8] ), .IN2(\r[21][8] ), .IN4(
        \r[23][8] ), .S0(n2046), .S1(n2027), .Q(n1646) );
  MUX41X1 U2131 ( .IN1(\r[16][8] ), .IN3(\r[18][8] ), .IN2(\r[17][8] ), .IN4(
        \r[19][8] ), .S0(n2046), .S1(n2027), .Q(n1647) );
  MUX41X1 U2132 ( .IN1(n1647), .IN3(n1645), .IN2(n1646), .IN4(n1644), .S0(N19),
        .S1(n2054), .Q(n1648) );
  MUX41X1 U2133 ( .IN1(\r[12][8] ), .IN3(\r[14][8] ), .IN2(\r[13][8] ), .IN4(
        \r[15][8] ), .S0(n2046), .S1(n2027), .Q(n1649) );
  MUX41X1 U2134 ( .IN1(\r[8][8] ), .IN3(\r[10][8] ), .IN2(\r[9][8] ), .IN4(
        \r[11][8] ), .S0(n2046), .S1(n2028), .Q(n1650) );
  MUX41X1 U2135 ( .IN1(\r[4][8] ), .IN3(\r[6][8] ), .IN2(\r[5][8] ), .IN4(
        \r[7][8] ), .S0(n2046), .S1(n2028), .Q(n1651) );
  MUX41X1 U2136 ( .IN1(n1652), .IN3(n1650), .IN2(n1651), .IN4(n1649), .S0(N19),
        .S1(n2054), .Q(n1653) );
  MUX21X1 U2137 ( .IN1(n1653), .IN2(n1648), .S(N20), .Q(rd_dataB[8]) );
  MUX41X1 U2138 ( .IN1(\r[28][9] ), .IN3(\r[30][9] ), .IN2(\r[29][9] ), .IN4(
        \r[31][9] ), .S0(n2046), .S1(n2028), .Q(n1654) );
  MUX41X1 U2139 ( .IN1(\r[24][9] ), .IN3(\r[26][9] ), .IN2(\r[25][9] ), .IN4(
        \r[27][9] ), .S0(n2046), .S1(n2028), .Q(n1655) );
  MUX41X1 U2140 ( .IN1(\r[20][9] ), .IN3(\r[22][9] ), .IN2(\r[21][9] ), .IN4(
        \r[23][9] ), .S0(n2046), .S1(n2028), .Q(n1656) );
  MUX41X1 U2141 ( .IN1(\r[16][9] ), .IN3(\r[18][9] ), .IN2(\r[17][9] ), .IN4(
        \r[19][9] ), .S0(n2046), .S1(n2028), .Q(n1657) );
  MUX41X1 U2142 ( .IN1(n1657), .IN3(n1655), .IN2(n1656), .IN4(n1654), .S0(N19),
        .S1(n2054), .Q(n1658) );
  MUX41X1 U2143 ( .IN1(\r[12][9] ), .IN3(\r[14][9] ), .IN2(\r[13][9] ), .IN4(
        \r[15][9] ), .S0(n2046), .S1(n2028), .Q(n1659) );
  MUX41X1 U2144 ( .IN1(\r[8][9] ), .IN3(\r[10][9] ), .IN2(\r[9][9] ), .IN4(
        \r[11][9] ), .S0(n2046), .S1(n2028), .Q(n1660) );
  MUX41X1 U2145 ( .IN1(\r[4][9] ), .IN3(\r[6][9] ), .IN2(\r[5][9] ), .IN4(
        \r[7][9] ), .S0(n2046), .S1(n2028), .Q(n1661) );
  MUX41X1 U2146 ( .IN1(n1662), .IN3(n1660), .IN2(n1661), .IN4(n1659), .S0(N19),
        .S1(n2054), .Q(n1663) );
  MUX21X1 U2147 ( .IN1(n1663), .IN2(n1658), .S(N20), .Q(rd_dataB[9]) );
  MUX41X1 U2148 ( .IN1(\r[28][10] ), .IN3(\r[30][10] ), .IN2(\r[29][10] ),
        .IN4(\r[31][10] ), .S0(n2046), .S1(n2028), .Q(n1664) );
  MUX41X1 U2149 ( .IN1(\r[24][10] ), .IN3(\r[26][10] ), .IN2(\r[25][10] ),
        .IN4(\r[27][10] ), .S0(n2046), .S1(n2028), .Q(n1665) );
  MUX41X1 U2150 ( .IN1(\r[20][10] ), .IN3(\r[22][10] ), .IN2(\r[21][10] ),
        .IN4(\r[23][10] ), .S0(n2046), .S1(n2028), .Q(n1666) );
  MUX41X1 U2151 ( .IN1(\r[16][10] ), .IN3(\r[18][10] ), .IN2(\r[17][10] ),
        .IN4(\r[19][10] ), .S0(n2046), .S1(n2029), .Q(n1667) );
  MUX41X1 U2152 ( .IN1(n1667), .IN3(n1665), .IN2(n1666), .IN4(n1664), .S0(N19),
        .S1(n2054), .Q(n1668) );
  MUX41X1 U2153 ( .IN1(\r[12][10] ), .IN3(\r[14][10] ), .IN2(\r[13][10] ),
        .IN4(\r[15][10] ), .S0(n2046), .S1(n2029), .Q(n1669) );
  MUX41X1 U2154 ( .IN1(\r[8][10] ), .IN3(\r[10][10] ), .IN2(\r[9][10] ), .IN4(
        \r[11][10] ), .S0(n2046), .S1(n2029), .Q(n1670) );
  MUX41X1 U2155 ( .IN1(\r[4][10] ), .IN3(\r[6][10] ), .IN2(\r[5][10] ), .IN4(
        \r[7][10] ), .S0(n2047), .S1(n2029), .Q(n1671) );
  MUX41X1 U2156 ( .IN1(n1672), .IN3(n1670), .IN2(n1671), .IN4(n1669), .S0(N19),
        .S1(n2054), .Q(n1673) );
  MUX21X1 U2157 ( .IN1(n1673), .IN2(n1668), .S(N20), .Q(rd_dataB[10]) );
  MUX41X1 U2158 ( .IN1(\r[28][11] ), .IN3(\r[30][11] ), .IN2(\r[29][11] ),
        .IN4(\r[31][11] ), .S0(n2047), .S1(n2029), .Q(n1674) );
  MUX41X1 U2159 ( .IN1(\r[24][11] ), .IN3(\r[26][11] ), .IN2(\r[25][11] ),
        .IN4(\r[27][11] ), .S0(n2047), .S1(n2029), .Q(n1675) );
  MUX41X1 U2160 ( .IN1(\r[20][11] ), .IN3(\r[22][11] ), .IN2(\r[21][11] ),
        .IN4(\r[23][11] ), .S0(n2047), .S1(n2029), .Q(n1676) );
  MUX41X1 U2161 ( .IN1(\r[16][11] ), .IN3(\r[18][11] ), .IN2(\r[17][11] ),
        .IN4(\r[19][11] ), .S0(n2047), .S1(n2029), .Q(n1677) );
  MUX41X1 U2162 ( .IN1(n1677), .IN3(n1675), .IN2(n1676), .IN4(n1674), .S0(N19),
        .S1(n2054), .Q(n1678) );
  MUX41X1 U2163 ( .IN1(\r[12][11] ), .IN3(\r[14][11] ), .IN2(\r[13][11] ),
        .IN4(\r[15][11] ), .S0(n2047), .S1(n2029), .Q(n1679) );
  MUX41X1 U2164 ( .IN1(\r[8][11] ), .IN3(\r[10][11] ), .IN2(\r[9][11] ), .IN4(
        \r[11][11] ), .S0(n2047), .S1(n2029), .Q(n1680) );
  MUX41X1 U2165 ( .IN1(\r[4][11] ), .IN3(\r[6][11] ), .IN2(\r[5][11] ), .IN4(
        \r[7][11] ), .S0(n2047), .S1(n2029), .Q(n1681) );
  MUX41X1 U2166 ( .IN1(n1682), .IN3(n1680), .IN2(n1681), .IN4(n1679), .S0(N19),
        .S1(n2054), .Q(n1683) );
  MUX21X1 U2167 ( .IN1(n1683), .IN2(n1678), .S(N20), .Q(rd_dataB[11]) );
  MUX41X1 U2168 ( .IN1(\r[28][12] ), .IN3(\r[30][12] ), .IN2(\r[29][12] ),
        .IN4(\r[31][12] ), .S0(n2047), .S1(n2030), .Q(n1684) );
  MUX41X1 U2169 ( .IN1(\r[24][12] ), .IN3(\r[26][12] ), .IN2(\r[25][12] ),
        .IN4(\r[27][12] ), .S0(n2047), .S1(n2030), .Q(n1685) );
  MUX41X1 U2170 ( .IN1(\r[20][12] ), .IN3(\r[22][12] ), .IN2(\r[21][12] ),
        .IN4(\r[23][12] ), .S0(n2047), .S1(n2030), .Q(n1686) );
  MUX41X1 U2171 ( .IN1(\r[16][12] ), .IN3(\r[18][12] ), .IN2(\r[17][12] ),
        .IN4(\r[19][12] ), .S0(n2047), .S1(n2030), .Q(n1687) );
  MUX41X1 U2172 ( .IN1(n1687), .IN3(n1685), .IN2(n1686), .IN4(n1684), .S0(N19),
        .S1(n2053), .Q(n1688) );
  MUX41X1 U2173 ( .IN1(\r[12][12] ), .IN3(\r[14][12] ), .IN2(\r[13][12] ),
        .IN4(\r[15][12] ), .S0(n2047), .S1(n2030), .Q(n1689) );
  MUX41X1 U2174 ( .IN1(\r[8][12] ), .IN3(\r[10][12] ), .IN2(\r[9][12] ), .IN4(
        \r[11][12] ), .S0(n2047), .S1(n2030), .Q(n1690) );
  MUX41X1 U2175 ( .IN1(\r[4][12] ), .IN3(\r[6][12] ), .IN2(\r[5][12] ), .IN4(
        \r[7][12] ), .S0(n2047), .S1(n2030), .Q(n1691) );
  MUX41X1 U2176 ( .IN1(n1692), .IN3(n1690), .IN2(n1691), .IN4(n1689), .S0(N19),
        .S1(n2053), .Q(n1693) );
  MUX21X1 U2177 ( .IN1(n1693), .IN2(n1688), .S(N20), .Q(rd_dataB[12]) );
  MUX41X1 U2178 ( .IN1(\r[28][13] ), .IN3(\r[30][13] ), .IN2(\r[29][13] ),
        .IN4(\r[31][13] ), .S0(n2047), .S1(n2030), .Q(n1694) );
  MUX41X1 U2179 ( .IN1(\r[24][13] ), .IN3(\r[26][13] ), .IN2(\r[25][13] ),
        .IN4(\r[27][13] ), .S0(n2047), .S1(n2030), .Q(n1695) );
  MUX41X1 U2180 ( .IN1(\r[20][13] ), .IN3(\r[22][13] ), .IN2(\r[21][13] ),
        .IN4(\r[23][13] ), .S0(n2047), .S1(n2030), .Q(n1696) );
  MUX41X1 U2181 ( .IN1(\r[16][13] ), .IN3(\r[18][13] ), .IN2(\r[17][13] ),
        .IN4(\r[19][13] ), .S0(n2047), .S1(n2030), .Q(n1697) );
  MUX41X1 U2182 ( .IN1(n1697), .IN3(n1695), .IN2(n1696), .IN4(n1694), .S0(N19),
        .S1(n2053), .Q(n1698) );
  MUX41X1 U2183 ( .IN1(\r[12][13] ), .IN3(\r[14][13] ), .IN2(\r[13][13] ),
        .IN4(\r[15][13] ), .S0(n2047), .S1(n2030), .Q(n1699) );
  MUX41X1 U2184 ( .IN1(\r[8][13] ), .IN3(\r[10][13] ), .IN2(\r[9][13] ), .IN4(
        \r[11][13] ), .S0(n2047), .S1(n2031), .Q(n1700) );
  MUX41X1 U2185 ( .IN1(\r[4][13] ), .IN3(\r[6][13] ), .IN2(\r[5][13] ), .IN4(
        \r[7][13] ), .S0(n2048), .S1(n2031), .Q(n1701) );
  MUX41X1 U2186 ( .IN1(n1702), .IN3(n1700), .IN2(n1701), .IN4(n1699), .S0(N19),
        .S1(n2053), .Q(n1703) );
  MUX21X1 U2187 ( .IN1(n1703), .IN2(n1698), .S(N20), .Q(rd_dataB[13]) );
  MUX41X1 U2188 ( .IN1(\r[28][14] ), .IN3(\r[30][14] ), .IN2(\r[29][14] ),
        .IN4(\r[31][14] ), .S0(n2047), .S1(n2031), .Q(n1704) );
  MUX41X1 U2189 ( .IN1(\r[24][14] ), .IN3(\r[26][14] ), .IN2(\r[25][14] ),
        .IN4(\r[27][14] ), .S0(n2048), .S1(n2031), .Q(n1705) );
  MUX41X1 U2190 ( .IN1(\r[20][14] ), .IN3(\r[22][14] ), .IN2(\r[21][14] ),
        .IN4(\r[23][14] ), .S0(n2048), .S1(n2031), .Q(n1706) );
  MUX41X1 U2191 ( .IN1(\r[16][14] ), .IN3(\r[18][14] ), .IN2(\r[17][14] ),
        .IN4(\r[19][14] ), .S0(n2048), .S1(n2031), .Q(n1707) );
  MUX41X1 U2192 ( .IN1(n1707), .IN3(n1705), .IN2(n1706), .IN4(n1704), .S0(N19),
        .S1(n2053), .Q(n1708) );
  MUX41X1 U2193 ( .IN1(\r[12][14] ), .IN3(\r[14][14] ), .IN2(\r[13][14] ),
        .IN4(\r[15][14] ), .S0(n2048), .S1(n2031), .Q(n1709) );
  MUX41X1 U2194 ( .IN1(\r[8][14] ), .IN3(\r[10][14] ), .IN2(\r[9][14] ), .IN4(
        \r[11][14] ), .S0(n2048), .S1(n2031), .Q(n1710) );
  MUX41X1 U2195 ( .IN1(\r[4][14] ), .IN3(\r[6][14] ), .IN2(\r[5][14] ), .IN4(
        \r[7][14] ), .S0(n2048), .S1(n2031), .Q(n1711) );
  MUX41X1 U2196 ( .IN1(n1712), .IN3(n1710), .IN2(n1711), .IN4(n1709), .S0(N19),
        .S1(n2053), .Q(n1713) );
  MUX21X1 U2197 ( .IN1(n1713), .IN2(n1708), .S(N20), .Q(rd_dataB[14]) );
  MUX41X1 U2198 ( .IN1(\r[28][15] ), .IN3(\r[30][15] ), .IN2(\r[29][15] ),
        .IN4(\r[31][15] ), .S0(n2048), .S1(n2031), .Q(n1714) );
  MUX41X1 U2199 ( .IN1(\r[24][15] ), .IN3(\r[26][15] ), .IN2(\r[25][15] ),
        .IN4(\r[27][15] ), .S0(n2048), .S1(n2031), .Q(n1715) );
  MUX41X1 U2200 ( .IN1(\r[20][15] ), .IN3(\r[22][15] ), .IN2(\r[21][15] ),
        .IN4(\r[23][15] ), .S0(n2048), .S1(n2031), .Q(n1716) );
  MUX41X1 U2201 ( .IN1(\r[16][15] ), .IN3(\r[18][15] ), .IN2(\r[17][15] ),
        .IN4(\r[19][15] ), .S0(n2048), .S1(n2032), .Q(n1717) );
  MUX41X1 U2202 ( .IN1(n1717), .IN3(n1715), .IN2(n1716), .IN4(n1714), .S0(N19),
        .S1(n2053), .Q(n1718) );
  MUX41X1 U2203 ( .IN1(\r[12][15] ), .IN3(\r[14][15] ), .IN2(\r[13][15] ),
        .IN4(\r[15][15] ), .S0(n2048), .S1(n2032), .Q(n1719) );
  MUX41X1 U2204 ( .IN1(\r[8][15] ), .IN3(\r[10][15] ), .IN2(\r[9][15] ), .IN4(
        \r[11][15] ), .S0(n2048), .S1(n2032), .Q(n1720) );
  MUX41X1 U2205 ( .IN1(\r[4][15] ), .IN3(\r[6][15] ), .IN2(\r[5][15] ), .IN4(
        \r[7][15] ), .S0(n2048), .S1(n2032), .Q(n1721) );
  MUX41X1 U2206 ( .IN1(n1722), .IN3(n1720), .IN2(n1721), .IN4(n1719), .S0(N19),
        .S1(n2053), .Q(n1723) );
  MUX21X1 U2207 ( .IN1(n1723), .IN2(n1718), .S(N20), .Q(rd_dataB[15]) );
  MUX41X1 U2208 ( .IN1(\r[28][16] ), .IN3(\r[30][16] ), .IN2(\r[29][16] ),
        .IN4(\r[31][16] ), .S0(n2048), .S1(n2032), .Q(n1724) );
  MUX41X1 U2209 ( .IN1(\r[24][16] ), .IN3(\r[26][16] ), .IN2(\r[25][16] ),
        .IN4(\r[27][16] ), .S0(n2048), .S1(n2032), .Q(n1725) );
  MUX41X1 U2210 ( .IN1(\r[20][16] ), .IN3(\r[22][16] ), .IN2(\r[21][16] ),
        .IN4(\r[23][16] ), .S0(n2048), .S1(n2032), .Q(n1726) );
  MUX41X1 U2211 ( .IN1(\r[16][16] ), .IN3(\r[18][16] ), .IN2(\r[17][16] ),
        .IN4(\r[19][16] ), .S0(n2049), .S1(n2032), .Q(n1727) );
  MUX41X1 U2212 ( .IN1(n1727), .IN3(n1725), .IN2(n1726), .IN4(n1724), .S0(N19),
        .S1(n2053), .Q(n1728) );
  MUX41X1 U2213 ( .IN1(\r[12][16] ), .IN3(\r[14][16] ), .IN2(\r[13][16] ),
        .IN4(\r[15][16] ), .S0(n2048), .S1(n2032), .Q(n1729) );
  MUX41X1 U2214 ( .IN1(\r[8][16] ), .IN3(\r[10][16] ), .IN2(\r[9][16] ), .IN4(
        \r[11][16] ), .S0(n2049), .S1(n2032), .Q(n1730) );
  MUX41X1 U2215 ( .IN1(\r[4][16] ), .IN3(\r[6][16] ), .IN2(\r[5][16] ), .IN4(
        \r[7][16] ), .S0(n2048), .S1(n2032), .Q(n1731) );
  MUX41X1 U2216 ( .IN1(n1732), .IN3(n1730), .IN2(n1731), .IN4(n1729), .S0(N19),
        .S1(n2053), .Q(n1733) );
  MUX21X1 U2217 ( .IN1(n1733), .IN2(n1728), .S(N20), .Q(rd_dataB[16]) );
  MUX41X1 U2218 ( .IN1(\r[28][17] ), .IN3(\r[30][17] ), .IN2(\r[29][17] ),
        .IN4(\r[31][17] ), .S0(n2048), .S1(n2032), .Q(n1734) );
  MUX41X1 U2219 ( .IN1(\r[24][17] ), .IN3(\r[26][17] ), .IN2(\r[25][17] ),
        .IN4(\r[27][17] ), .S0(n2049), .S1(n2033), .Q(n1735) );
  MUX41X1 U2220 ( .IN1(\r[20][17] ), .IN3(\r[22][17] ), .IN2(\r[21][17] ),
        .IN4(\r[23][17] ), .S0(n2049), .S1(n2033), .Q(n1736) );
  MUX41X1 U2221 ( .IN1(\r[16][17] ), .IN3(\r[18][17] ), .IN2(\r[17][17] ),
        .IN4(\r[19][17] ), .S0(n2048), .S1(n2033), .Q(n1737) );
  MUX41X1 U2222 ( .IN1(n1737), .IN3(n1735), .IN2(n1736), .IN4(n1734), .S0(N19),
        .S1(n2053), .Q(n1738) );
  MUX41X1 U2223 ( .IN1(\r[12][17] ), .IN3(\r[14][17] ), .IN2(\r[13][17] ),
        .IN4(\r[15][17] ), .S0(n2049), .S1(n2033), .Q(n1739) );
  MUX41X1 U2224 ( .IN1(\r[8][17] ), .IN3(\r[10][17] ), .IN2(\r[9][17] ), .IN4(
        \r[11][17] ), .S0(n2049), .S1(n2033), .Q(n1740) );
  MUX41X1 U2225 ( .IN1(\r[4][17] ), .IN3(\r[6][17] ), .IN2(\r[5][17] ), .IN4(
        \r[7][17] ), .S0(n2048), .S1(n2033), .Q(n1741) );
  MUX41X1 U2226 ( .IN1(n1742), .IN3(n1740), .IN2(n1741), .IN4(n1739), .S0(N19),
        .S1(n2053), .Q(n1743) );
  MUX21X1 U2227 ( .IN1(n1743), .IN2(n1738), .S(N20), .Q(rd_dataB[17]) );
  MUX41X1 U2228 ( .IN1(\r[28][18] ), .IN3(\r[30][18] ), .IN2(\r[29][18] ),
        .IN4(\r[31][18] ), .S0(n2049), .S1(n2033), .Q(n1744) );
  MUX41X1 U2229 ( .IN1(\r[24][18] ), .IN3(\r[26][18] ), .IN2(\r[25][18] ),
        .IN4(\r[27][18] ), .S0(n2046), .S1(n2033), .Q(n1745) );
  MUX41X1 U2230 ( .IN1(\r[20][18] ), .IN3(\r[22][18] ), .IN2(\r[21][18] ),
        .IN4(\r[23][18] ), .S0(n2039), .S1(n2033), .Q(n1746) );
  MUX41X1 U2231 ( .IN1(\r[16][18] ), .IN3(\r[18][18] ), .IN2(\r[17][18] ),
        .IN4(\r[19][18] ), .S0(n2039), .S1(n2033), .Q(n1747) );
  MUX41X1 U2232 ( .IN1(n1747), .IN3(n1745), .IN2(n1746), .IN4(n1744), .S0(N19),
        .S1(n2052), .Q(n1748) );
  MUX41X1 U2233 ( .IN1(\r[12][18] ), .IN3(\r[14][18] ), .IN2(\r[13][18] ),
        .IN4(\r[15][18] ), .S0(n2039), .S1(n2033), .Q(n1749) );
  MUX41X1 U2234 ( .IN1(\r[8][18] ), .IN3(\r[10][18] ), .IN2(\r[9][18] ), .IN4(
        \r[11][18] ), .S0(n2039), .S1(n2033), .Q(n1750) );
  MUX41X1 U2235 ( .IN1(\r[4][18] ), .IN3(\r[6][18] ), .IN2(\r[5][18] ), .IN4(
        \r[7][18] ), .S0(n2039), .S1(n2034), .Q(n1751) );
  MUX41X1 U2236 ( .IN1(n1752), .IN3(n1750), .IN2(n1751), .IN4(n1749), .S0(N19),
        .S1(n2052), .Q(n1753) );
  MUX21X1 U2237 ( .IN1(n1753), .IN2(n1748), .S(N20), .Q(rd_dataB[18]) );
  MUX41X1 U2238 ( .IN1(\r[28][19] ), .IN3(\r[30][19] ), .IN2(\r[29][19] ),
        .IN4(\r[31][19] ), .S0(n2039), .S1(n2034), .Q(n1754) );
  MUX41X1 U2239 ( .IN1(\r[24][19] ), .IN3(\r[26][19] ), .IN2(\r[25][19] ),
        .IN4(\r[27][19] ), .S0(n2039), .S1(n2034), .Q(n1755) );
  MUX41X1 U2240 ( .IN1(\r[20][19] ), .IN3(\r[22][19] ), .IN2(\r[21][19] ),
        .IN4(\r[23][19] ), .S0(n2039), .S1(n2034), .Q(n1756) );
  MUX41X1 U2241 ( .IN1(\r[16][19] ), .IN3(\r[18][19] ), .IN2(\r[17][19] ),
        .IN4(\r[19][19] ), .S0(n2039), .S1(n2034), .Q(n1757) );
  MUX41X1 U2242 ( .IN1(n1757), .IN3(n1755), .IN2(n1756), .IN4(n1754), .S0(N19),
        .S1(n2052), .Q(n1758) );
  MUX41X1 U2243 ( .IN1(\r[12][19] ), .IN3(\r[14][19] ), .IN2(\r[13][19] ),
        .IN4(\r[15][19] ), .S0(n2039), .S1(n2034), .Q(n1759) );
  MUX41X1 U2244 ( .IN1(\r[8][19] ), .IN3(\r[10][19] ), .IN2(\r[9][19] ), .IN4(
        \r[11][19] ), .S0(n2039), .S1(n2034), .Q(n1760) );
  MUX41X1 U2245 ( .IN1(\r[4][19] ), .IN3(\r[6][19] ), .IN2(\r[5][19] ), .IN4(
        \r[7][19] ), .S0(n2039), .S1(n2034), .Q(n1761) );
  MUX41X1 U2246 ( .IN1(n1762), .IN3(n1760), .IN2(n1761), .IN4(n1759), .S0(N19),
        .S1(n2052), .Q(n1763) );
  MUX21X1 U2247 ( .IN1(n1763), .IN2(n1758), .S(N20), .Q(rd_dataB[19]) );
  MUX41X1 U2248 ( .IN1(\r[28][20] ), .IN3(\r[30][20] ), .IN2(\r[29][20] ),
        .IN4(\r[31][20] ), .S0(n2039), .S1(n2034), .Q(n1764) );
  MUX41X1 U2249 ( .IN1(\r[24][20] ), .IN3(\r[26][20] ), .IN2(\r[25][20] ),
        .IN4(\r[27][20] ), .S0(n2039), .S1(n2034), .Q(n1765) );
  MUX41X1 U2250 ( .IN1(\r[20][20] ), .IN3(\r[22][20] ), .IN2(\r[21][20] ),
        .IN4(\r[23][20] ), .S0(n2039), .S1(n2034), .Q(n1766) );
  MUX41X1 U2251 ( .IN1(\r[16][20] ), .IN3(\r[18][20] ), .IN2(\r[17][20] ),
        .IN4(\r[19][20] ), .S0(n2039), .S1(n2029), .Q(n1767) );
  MUX41X1 U2252 ( .IN1(n1767), .IN3(n1765), .IN2(n1766), .IN4(n1764), .S0(N19),
        .S1(n2052), .Q(n1768) );
  MUX41X1 U2253 ( .IN1(\r[12][20] ), .IN3(\r[14][20] ), .IN2(\r[13][20] ),
        .IN4(\r[15][20] ), .S0(n2041), .S1(n2020), .Q(n1769) );
  MUX41X1 U2254 ( .IN1(\r[8][20] ), .IN3(\r[10][20] ), .IN2(\r[9][20] ), .IN4(
        \r[11][20] ), .S0(n2039), .S1(n2017), .Q(n1770) );
  MUX41X1 U2255 ( .IN1(\r[4][20] ), .IN3(\r[6][20] ), .IN2(\r[5][20] ), .IN4(
        \r[7][20] ), .S0(n2040), .S1(n2017), .Q(n1771) );
  MUX41X1 U2256 ( .IN1(n1772), .IN3(n1770), .IN2(n1771), .IN4(n1769), .S0(N19),
        .S1(n2052), .Q(n1773) );
  MUX21X1 U2257 ( .IN1(n1773), .IN2(n1768), .S(N20), .Q(rd_dataB[20]) );
  MUX41X1 U2258 ( .IN1(\r[28][21] ), .IN3(\r[30][21] ), .IN2(\r[29][21] ),
        .IN4(\r[31][21] ), .S0(n2040), .S1(n2017), .Q(n1774) );
  MUX41X1 U2259 ( .IN1(\r[24][21] ), .IN3(\r[26][21] ), .IN2(\r[25][21] ),
        .IN4(\r[27][21] ), .S0(n2040), .S1(n2017), .Q(n1775) );
  MUX41X1 U2260 ( .IN1(\r[20][21] ), .IN3(\r[22][21] ), .IN2(\r[21][21] ),
        .IN4(\r[23][21] ), .S0(n2040), .S1(n2017), .Q(n1776) );
  MUX41X1 U2261 ( .IN1(\r[16][21] ), .IN3(\r[18][21] ), .IN2(\r[17][21] ),
        .IN4(\r[19][21] ), .S0(n2040), .S1(n2017), .Q(n1777) );
  MUX41X1 U2262 ( .IN1(n1777), .IN3(n1775), .IN2(n1776), .IN4(n1774), .S0(N19),
        .S1(n2052), .Q(n1778) );
  MUX41X1 U2263 ( .IN1(\r[12][21] ), .IN3(\r[14][21] ), .IN2(\r[13][21] ),
        .IN4(\r[15][21] ), .S0(n2040), .S1(n2017), .Q(n1779) );
  MUX41X1 U2264 ( .IN1(\r[8][21] ), .IN3(\r[10][21] ), .IN2(\r[9][21] ), .IN4(
        \r[11][21] ), .S0(n2040), .S1(n2018), .Q(n1780) );
  MUX41X1 U2265 ( .IN1(\r[4][21] ), .IN3(\r[6][21] ), .IN2(\r[5][21] ), .IN4(
        \r[7][21] ), .S0(n2040), .S1(n2018), .Q(n1781) );
  MUX41X1 U2266 ( .IN1(n1782), .IN3(n1780), .IN2(n1781), .IN4(n1779), .S0(N19),
        .S1(n2052), .Q(n1783) );
  MUX21X1 U2267 ( .IN1(n1783), .IN2(n1778), .S(N20), .Q(rd_dataB[21]) );
  MUX41X1 U2268 ( .IN1(\r[28][22] ), .IN3(\r[30][22] ), .IN2(\r[29][22] ),
        .IN4(\r[31][22] ), .S0(n2040), .S1(n2018), .Q(n1784) );
  MUX41X1 U2269 ( .IN1(\r[24][22] ), .IN3(\r[26][22] ), .IN2(\r[25][22] ),
        .IN4(\r[27][22] ), .S0(n2040), .S1(n2018), .Q(n1785) );
  MUX41X1 U2270 ( .IN1(\r[20][22] ), .IN3(\r[22][22] ), .IN2(\r[21][22] ),
        .IN4(\r[23][22] ), .S0(n2040), .S1(n2018), .Q(n1786) );
  MUX41X1 U2271 ( .IN1(\r[16][22] ), .IN3(\r[18][22] ), .IN2(\r[17][22] ),
        .IN4(\r[19][22] ), .S0(n2040), .S1(n2018), .Q(n1787) );
  MUX41X1 U2272 ( .IN1(n1787), .IN3(n1785), .IN2(n1786), .IN4(n1784), .S0(N19),
        .S1(n2052), .Q(n1788) );
  MUX41X1 U2273 ( .IN1(\r[12][22] ), .IN3(\r[14][22] ), .IN2(\r[13][22] ),
        .IN4(\r[15][22] ), .S0(n2040), .S1(n2018), .Q(n1789) );
  MUX41X1 U2274 ( .IN1(\r[8][22] ), .IN3(\r[10][22] ), .IN2(\r[9][22] ), .IN4(
        \r[11][22] ), .S0(n2040), .S1(n2018), .Q(n1790) );
  MUX41X1 U2275 ( .IN1(\r[4][22] ), .IN3(\r[6][22] ), .IN2(\r[5][22] ), .IN4(
        \r[7][22] ), .S0(n2040), .S1(n2018), .Q(n1791) );
  MUX41X1 U2276 ( .IN1(n1792), .IN3(n1790), .IN2(n1791), .IN4(n1789), .S0(N19),
        .S1(n2052), .Q(n1793) );
  MUX21X1 U2277 ( .IN1(n1793), .IN2(n1788), .S(N20), .Q(rd_dataB[22]) );
  MUX41X1 U2278 ( .IN1(\r[28][23] ), .IN3(\r[30][23] ), .IN2(\r[29][23] ),
        .IN4(\r[31][23] ), .S0(n2040), .S1(n2018), .Q(n1794) );
  MUX41X1 U2279 ( .IN1(\r[24][23] ), .IN3(\r[26][23] ), .IN2(\r[25][23] ),
        .IN4(\r[27][23] ), .S0(n2040), .S1(n2018), .Q(n1795) );
  MUX41X1 U2280 ( .IN1(\r[20][23] ), .IN3(\r[22][23] ), .IN2(\r[21][23] ),
        .IN4(\r[23][23] ), .S0(n2040), .S1(n2018), .Q(n1796) );
  MUX41X1 U2281 ( .IN1(\r[16][23] ), .IN3(\r[18][23] ), .IN2(\r[17][23] ),
        .IN4(\r[19][23] ), .S0(n2040), .S1(n2019), .Q(n1797) );
  MUX41X1 U2282 ( .IN1(n1797), .IN3(n1795), .IN2(n1796), .IN4(n1794), .S0(N19),
        .S1(n2052), .Q(n1798) );
  MUX41X1 U2283 ( .IN1(\r[12][23] ), .IN3(\r[14][23] ), .IN2(\r[13][23] ),
        .IN4(\r[15][23] ), .S0(n2040), .S1(n2019), .Q(n1799) );
  MUX41X1 U2284 ( .IN1(\r[8][23] ), .IN3(\r[10][23] ), .IN2(\r[9][23] ), .IN4(
        \r[11][23] ), .S0(n2040), .S1(n2019), .Q(n1800) );
  MUX41X1 U2285 ( .IN1(\r[4][23] ), .IN3(\r[6][23] ), .IN2(\r[5][23] ), .IN4(
        \r[7][23] ), .S0(n2040), .S1(n2019), .Q(n1801) );
  MUX41X1 U2286 ( .IN1(n1802), .IN3(n1800), .IN2(n1801), .IN4(n1799), .S0(N19),
        .S1(n2052), .Q(n1803) );
  MUX21X1 U2287 ( .IN1(n1803), .IN2(n1798), .S(N20), .Q(rd_dataB[23]) );
  MUX41X1 U2288 ( .IN1(\r[28][24] ), .IN3(\r[30][24] ), .IN2(\r[29][24] ),
        .IN4(\r[31][24] ), .S0(n2041), .S1(n2019), .Q(n1804) );
  MUX41X1 U2289 ( .IN1(\r[24][24] ), .IN3(\r[26][24] ), .IN2(\r[25][24] ),
        .IN4(\r[27][24] ), .S0(n2041), .S1(n2019), .Q(n1805) );
  MUX41X1 U2290 ( .IN1(\r[20][24] ), .IN3(\r[22][24] ), .IN2(\r[21][24] ),
        .IN4(\r[23][24] ), .S0(n2041), .S1(n2019), .Q(n1806) );
  MUX41X1 U2291 ( .IN1(\r[16][24] ), .IN3(\r[18][24] ), .IN2(\r[17][24] ),
        .IN4(\r[19][24] ), .S0(n2041), .S1(n2019), .Q(n1807) );
  MUX41X1 U2292 ( .IN1(n1807), .IN3(n1805), .IN2(n1806), .IN4(n1804), .S0(N19),
        .S1(N18), .Q(n1808) );
  MUX41X1 U2293 ( .IN1(\r[12][24] ), .IN3(\r[14][24] ), .IN2(\r[13][24] ),
        .IN4(\r[15][24] ), .S0(n2041), .S1(n2019), .Q(n1809) );
  MUX41X1 U2294 ( .IN1(\r[8][24] ), .IN3(\r[10][24] ), .IN2(\r[9][24] ), .IN4(
        \r[11][24] ), .S0(n2041), .S1(n2019), .Q(n1810) );
  MUX41X1 U2295 ( .IN1(\r[4][24] ), .IN3(\r[6][24] ), .IN2(\r[5][24] ), .IN4(
        \r[7][24] ), .S0(n2041), .S1(n2019), .Q(n1811) );
  MUX41X1 U2296 ( .IN1(n1812), .IN3(n1810), .IN2(n1811), .IN4(n1809), .S0(N19),
        .S1(N18), .Q(n1813) );
  MUX21X1 U2297 ( .IN1(n1813), .IN2(n1808), .S(N20), .Q(rd_dataB[24]) );
  MUX41X1 U2298 ( .IN1(\r[28][25] ), .IN3(\r[30][25] ), .IN2(\r[29][25] ),
        .IN4(\r[31][25] ), .S0(n2041), .S1(n2019), .Q(n1814) );
  MUX41X1 U2299 ( .IN1(\r[24][25] ), .IN3(\r[26][25] ), .IN2(\r[25][25] ),
        .IN4(\r[27][25] ), .S0(n2041), .S1(n2020), .Q(n1815) );
  MUX41X1 U2300 ( .IN1(\r[20][25] ), .IN3(\r[22][25] ), .IN2(\r[21][25] ),
        .IN4(\r[23][25] ), .S0(n2041), .S1(n2020), .Q(n1816) );
  MUX41X1 U2301 ( .IN1(\r[16][25] ), .IN3(\r[18][25] ), .IN2(\r[17][25] ),
        .IN4(\r[19][25] ), .S0(n2041), .S1(n2020), .Q(n1817) );
  MUX41X1 U2302 ( .IN1(n1817), .IN3(n1815), .IN2(n1816), .IN4(n1814), .S0(N19),
        .S1(N18), .Q(n1818) );
  MUX41X1 U2303 ( .IN1(\r[12][25] ), .IN3(\r[14][25] ), .IN2(\r[13][25] ),
        .IN4(\r[15][25] ), .S0(n2041), .S1(n2020), .Q(n1819) );
  MUX41X1 U2304 ( .IN1(\r[8][25] ), .IN3(\r[10][25] ), .IN2(\r[9][25] ), .IN4(
        \r[11][25] ), .S0(n2041), .S1(n2020), .Q(n1820) );
  MUX41X1 U2305 ( .IN1(\r[4][25] ), .IN3(\r[6][25] ), .IN2(\r[5][25] ), .IN4(
        \r[7][25] ), .S0(n2041), .S1(n2020), .Q(n1821) );
  MUX41X1 U2306 ( .IN1(n1822), .IN3(n1820), .IN2(n1821), .IN4(n1819), .S0(N19),
        .S1(N18), .Q(n1823) );
  MUX21X1 U2307 ( .IN1(n1823), .IN2(n1818), .S(N20), .Q(rd_dataB[25]) );
  MUX41X1 U2308 ( .IN1(\r[28][26] ), .IN3(\r[30][26] ), .IN2(\r[29][26] ),
        .IN4(\r[31][26] ), .S0(n2041), .S1(n2020), .Q(n1824) );
  MUX41X1 U2309 ( .IN1(\r[24][26] ), .IN3(\r[26][26] ), .IN2(\r[25][26] ),
        .IN4(\r[27][26] ), .S0(n2041), .S1(n2020), .Q(n1825) );
  MUX41X1 U2310 ( .IN1(\r[20][26] ), .IN3(\r[22][26] ), .IN2(\r[21][26] ),
        .IN4(\r[23][26] ), .S0(n2041), .S1(n2020), .Q(n1826) );
  MUX41X1 U2311 ( .IN1(\r[16][26] ), .IN3(\r[18][26] ), .IN2(\r[17][26] ),
        .IN4(\r[19][26] ), .S0(n2041), .S1(n2020), .Q(n1827) );
  MUX41X1 U2312 ( .IN1(n1827), .IN3(n1825), .IN2(n1826), .IN4(n1824), .S0(N19),
        .S1(N18), .Q(n1828) );
  MUX41X1 U2313 ( .IN1(\r[12][26] ), .IN3(\r[14][26] ), .IN2(\r[13][26] ),
        .IN4(\r[15][26] ), .S0(n2041), .S1(n2020), .Q(n1829) );
  MUX41X1 U2314 ( .IN1(\r[8][26] ), .IN3(\r[10][26] ), .IN2(\r[9][26] ), .IN4(
        \r[11][26] ), .S0(n2041), .S1(n2021), .Q(n1830) );
  MUX41X1 U2315 ( .IN1(\r[4][26] ), .IN3(\r[6][26] ), .IN2(\r[5][26] ), .IN4(
        \r[7][26] ), .S0(n2041), .S1(n2021), .Q(n1831) );
  MUX41X1 U2316 ( .IN1(n1832), .IN3(n1830), .IN2(n1831), .IN4(n1829), .S0(N19),
        .S1(N18), .Q(n1833) );
  MUX21X1 U2317 ( .IN1(n1833), .IN2(n1828), .S(N20), .Q(rd_dataB[26]) );
  MUX41X1 U2318 ( .IN1(\r[28][27] ), .IN3(\r[30][27] ), .IN2(\r[29][27] ),
        .IN4(\r[31][27] ), .S0(n2042), .S1(n2021), .Q(n1834) );
  MUX41X1 U2319 ( .IN1(\r[24][27] ), .IN3(\r[26][27] ), .IN2(\r[25][27] ),
        .IN4(\r[27][27] ), .S0(n2042), .S1(n2021), .Q(n1835) );
  MUX41X1 U2320 ( .IN1(\r[20][27] ), .IN3(\r[22][27] ), .IN2(\r[21][27] ),
        .IN4(\r[23][27] ), .S0(n2042), .S1(n2021), .Q(n1836) );
  MUX41X1 U2321 ( .IN1(\r[16][27] ), .IN3(\r[18][27] ), .IN2(\r[17][27] ),
        .IN4(\r[19][27] ), .S0(n2042), .S1(n2021), .Q(n1837) );
  MUX41X1 U2322 ( .IN1(n1837), .IN3(n1835), .IN2(n1836), .IN4(n1834), .S0(N19),
        .S1(N18), .Q(n1838) );
  MUX41X1 U2323 ( .IN1(\r[12][27] ), .IN3(\r[14][27] ), .IN2(\r[13][27] ),
        .IN4(\r[15][27] ), .S0(n2042), .S1(n2021), .Q(n1839) );
  MUX41X1 U2324 ( .IN1(\r[8][27] ), .IN3(\r[10][27] ), .IN2(\r[9][27] ), .IN4(
        \r[11][27] ), .S0(n2042), .S1(n2021), .Q(n1840) );
  MUX41X1 U2325 ( .IN1(\r[4][27] ), .IN3(\r[6][27] ), .IN2(\r[5][27] ), .IN4(
        \r[7][27] ), .S0(n2042), .S1(n2021), .Q(n1841) );
  MUX41X1 U2326 ( .IN1(n1842), .IN3(n1840), .IN2(n1841), .IN4(n1839), .S0(N19),
        .S1(N18), .Q(n1843) );
  MUX21X1 U2327 ( .IN1(n1843), .IN2(n1838), .S(N20), .Q(rd_dataB[27]) );
  MUX41X1 U2328 ( .IN1(\r[28][28] ), .IN3(\r[30][28] ), .IN2(\r[29][28] ),
        .IN4(\r[31][28] ), .S0(n2042), .S1(n2021), .Q(n1844) );
  MUX41X1 U2329 ( .IN1(\r[24][28] ), .IN3(\r[26][28] ), .IN2(\r[25][28] ),
        .IN4(\r[27][28] ), .S0(n2042), .S1(n2021), .Q(n1845) );
  MUX41X1 U2330 ( .IN1(\r[20][28] ), .IN3(\r[22][28] ), .IN2(\r[21][28] ),
        .IN4(\r[23][28] ), .S0(n2042), .S1(n2021), .Q(n1846) );
  MUX41X1 U2331 ( .IN1(\r[16][28] ), .IN3(\r[18][28] ), .IN2(\r[17][28] ),
        .IN4(\r[19][28] ), .S0(n2042), .S1(n2022), .Q(n1847) );
  MUX41X1 U2332 ( .IN1(n1847), .IN3(n1845), .IN2(n1846), .IN4(n1844), .S0(N19),
        .S1(N18), .Q(n1848) );
  MUX41X1 U2333 ( .IN1(\r[12][28] ), .IN3(\r[14][28] ), .IN2(\r[13][28] ),
        .IN4(\r[15][28] ), .S0(n2042), .S1(n2022), .Q(n1849) );
  MUX41X1 U2334 ( .IN1(\r[8][28] ), .IN3(\r[10][28] ), .IN2(\r[9][28] ), .IN4(
        \r[11][28] ), .S0(n2042), .S1(n2022), .Q(n1850) );
  MUX41X1 U2335 ( .IN1(\r[4][28] ), .IN3(\r[6][28] ), .IN2(\r[5][28] ), .IN4(
        \r[7][28] ), .S0(n2042), .S1(n2022), .Q(n1851) );
  MUX41X1 U2336 ( .IN1(n1852), .IN3(n1850), .IN2(n1851), .IN4(n1849), .S0(N19),
        .S1(N18), .Q(n1853) );
  MUX21X1 U2337 ( .IN1(n1853), .IN2(n1848), .S(N20), .Q(rd_dataB[28]) );
  MUX41X1 U2338 ( .IN1(\r[28][29] ), .IN3(\r[30][29] ), .IN2(\r[29][29] ),
        .IN4(\r[31][29] ), .S0(n2042), .S1(n2022), .Q(n1854) );
  MUX41X1 U2339 ( .IN1(\r[24][29] ), .IN3(\r[26][29] ), .IN2(\r[25][29] ),
        .IN4(\r[27][29] ), .S0(n2042), .S1(n2022), .Q(n1855) );
  MUX41X1 U2340 ( .IN1(\r[20][29] ), .IN3(\r[22][29] ), .IN2(\r[21][29] ),
        .IN4(\r[23][29] ), .S0(n2042), .S1(n2022), .Q(n1856) );
  MUX41X1 U2341 ( .IN1(\r[16][29] ), .IN3(\r[18][29] ), .IN2(\r[17][29] ),
        .IN4(\r[19][29] ), .S0(n2042), .S1(n2022), .Q(n1857) );
  MUX41X1 U2342 ( .IN1(n1857), .IN3(n1855), .IN2(n1856), .IN4(n1854), .S0(N19),
        .S1(N18), .Q(n1858) );
  MUX41X1 U2343 ( .IN1(\r[12][29] ), .IN3(\r[14][29] ), .IN2(\r[13][29] ),
        .IN4(\r[15][29] ), .S0(n2042), .S1(n2022), .Q(n1859) );
  MUX41X1 U2344 ( .IN1(\r[8][29] ), .IN3(\r[10][29] ), .IN2(\r[9][29] ), .IN4(
        \r[11][29] ), .S0(n2042), .S1(n2022), .Q(n1860) );
  MUX41X1 U2345 ( .IN1(\r[4][29] ), .IN3(\r[6][29] ), .IN2(\r[5][29] ), .IN4(
        \r[7][29] ), .S0(n2042), .S1(n2022), .Q(n1861) );
  MUX41X1 U2346 ( .IN1(n1862), .IN3(n1860), .IN2(n1861), .IN4(n1859), .S0(N19),
        .S1(N18), .Q(n1863) );
  MUX21X1 U2347 ( .IN1(n1863), .IN2(n1858), .S(N20), .Q(rd_dataB[29]) );
  MUX41X1 U2348 ( .IN1(\r[28][30] ), .IN3(\r[30][30] ), .IN2(\r[29][30] ),
        .IN4(\r[31][30] ), .S0(n2042), .S1(n2022), .Q(n1864) );
  MUX41X1 U2349 ( .IN1(\r[24][30] ), .IN3(\r[26][30] ), .IN2(\r[25][30] ),
        .IN4(\r[27][30] ), .S0(n2043), .S1(n2023), .Q(n1865) );
  MUX41X1 U2350 ( .IN1(\r[20][30] ), .IN3(\r[22][30] ), .IN2(\r[21][30] ),
        .IN4(\r[23][30] ), .S0(n2043), .S1(n2023), .Q(n1866) );
  MUX41X1 U2351 ( .IN1(\r[16][30] ), .IN3(\r[18][30] ), .IN2(\r[17][30] ),
        .IN4(\r[19][30] ), .S0(n2043), .S1(n2023), .Q(n1867) );
  MUX41X1 U2352 ( .IN1(n1867), .IN3(n1865), .IN2(n1866), .IN4(n1864), .S0(N19),
        .S1(N18), .Q(n1868) );
  MUX41X1 U2353 ( .IN1(\r[12][30] ), .IN3(\r[14][30] ), .IN2(\r[13][30] ),
        .IN4(\r[15][30] ), .S0(n2043), .S1(n2023), .Q(n1869) );
  MUX41X1 U2354 ( .IN1(\r[8][30] ), .IN3(\r[10][30] ), .IN2(\r[9][30] ), .IN4(
        \r[11][30] ), .S0(n2043), .S1(n2023), .Q(n1870) );
  MUX41X1 U2355 ( .IN1(\r[4][30] ), .IN3(\r[6][30] ), .IN2(\r[5][30] ), .IN4(
        \r[7][30] ), .S0(n2043), .S1(n2023), .Q(n1871) );
  MUX41X1 U2356 ( .IN1(n1872), .IN3(n1870), .IN2(n1871), .IN4(n1869), .S0(N19),
        .S1(N18), .Q(n1873) );
  MUX21X1 U2357 ( .IN1(n1873), .IN2(n1868), .S(N20), .Q(rd_dataB[30]) );
  MUX41X1 U2358 ( .IN1(\r[28][31] ), .IN3(\r[30][31] ), .IN2(\r[29][31] ),
        .IN4(\r[31][31] ), .S0(n2043), .S1(n2023), .Q(n1874) );
  MUX41X1 U2359 ( .IN1(\r[24][31] ), .IN3(\r[26][31] ), .IN2(\r[25][31] ),
        .IN4(\r[27][31] ), .S0(n2043), .S1(n2023), .Q(n1875) );
  MUX41X1 U2360 ( .IN1(\r[20][31] ), .IN3(\r[22][31] ), .IN2(\r[21][31] ),
        .IN4(\r[23][31] ), .S0(n2043), .S1(n2023), .Q(n1876) );
  MUX41X1 U2361 ( .IN1(\r[16][31] ), .IN3(\r[18][31] ), .IN2(\r[17][31] ),
        .IN4(\r[19][31] ), .S0(n2043), .S1(n2023), .Q(n1877) );
  MUX41X1 U2362 ( .IN1(n1877), .IN3(n1875), .IN2(n1876), .IN4(n1874), .S0(N19),
        .S1(N18), .Q(n1878) );
  MUX41X1 U2363 ( .IN1(\r[12][31] ), .IN3(\r[14][31] ), .IN2(\r[13][31] ),
        .IN4(\r[15][31] ), .S0(n2043), .S1(n2023), .Q(n1879) );
  MUX41X1 U2364 ( .IN1(\r[8][31] ), .IN3(\r[10][31] ), .IN2(\r[9][31] ), .IN4(
        \r[11][31] ), .S0(n2043), .S1(n2023), .Q(n1880) );
  MUX41X1 U2365 ( .IN1(\r[4][31] ), .IN3(\r[6][31] ), .IN2(\r[5][31] ), .IN4(
        \r[7][31] ), .S0(n2043), .S1(N16), .Q(n1881) );
  MUX41X1 U2366 ( .IN1(n1882), .IN3(n1880), .IN2(n1881), .IN4(n1879), .S0(N19),
        .S1(N18), .Q(n1883) );
  MUX21X1 U2367 ( .IN1(n1883), .IN2(n1878), .S(N20), .Q(rd_dataB[31]) );
  MUX21X1 U2368 ( .IN1(n1884), .IN2(n1885), .S(n2017), .Q(n1887) );
  NAND3X0 U2369 ( .IN1(\r[3][31] ), .IN2(n2014), .IN3(n2039), .QN(n1886) );
  MUX21X1 U2370 ( .IN1(n1888), .IN2(n1889), .S(n2015), .Q(n1891) );
  NAND3X0 U2371 ( .IN1(\r[3][30] ), .IN2(n2014), .IN3(n2039), .QN(n1890) );
  MUX21X1 U2372 ( .IN1(n1892), .IN2(n1893), .S(n2015), .Q(n1895) );
  NAND3X0 U2373 ( .IN1(\r[3][29] ), .IN2(n2014), .IN3(n2039), .QN(n1894) );
  MUX21X1 U2374 ( .IN1(n1896), .IN2(n1897), .S(n2015), .Q(n1899) );
  NAND3X0 U2375 ( .IN1(\r[3][28] ), .IN2(n2014), .IN3(n2039), .QN(n1898) );
  MUX21X1 U2376 ( .IN1(n1900), .IN2(n1901), .S(n2015), .Q(n1903) );
  NAND3X0 U2377 ( .IN1(\r[3][27] ), .IN2(n2014), .IN3(n2038), .QN(n1902) );
  MUX21X1 U2378 ( .IN1(n1904), .IN2(n1905), .S(n2015), .Q(n1907) );
  NAND3X0 U2379 ( .IN1(\r[3][26] ), .IN2(n2014), .IN3(n2038), .QN(n1906) );
  MUX21X1 U2380 ( .IN1(n1908), .IN2(n1909), .S(n2015), .Q(n1911) );
  NAND3X0 U2381 ( .IN1(\r[3][25] ), .IN2(n2015), .IN3(n2038), .QN(n1910) );
  MUX21X1 U2382 ( .IN1(n1912), .IN2(n1913), .S(n2015), .Q(n1915) );
  NAND3X0 U2383 ( .IN1(\r[3][24] ), .IN2(n2014), .IN3(n2038), .QN(n1914) );
  MUX21X1 U2384 ( .IN1(n1916), .IN2(n1917), .S(n2015), .Q(n1919) );
  NAND3X0 U2385 ( .IN1(\r[3][23] ), .IN2(n2015), .IN3(n2038), .QN(n1918) );
  MUX21X1 U2386 ( .IN1(n1920), .IN2(n1921), .S(n2016), .Q(n1923) );
  NAND3X0 U2387 ( .IN1(\r[3][22] ), .IN2(n2015), .IN3(n2038), .QN(n1922) );
  MUX21X1 U2388 ( .IN1(n1924), .IN2(n1925), .S(n2016), .Q(n1927) );
  NAND3X0 U2389 ( .IN1(\r[3][21] ), .IN2(n2015), .IN3(n2038), .QN(n1926) );
  MUX21X1 U2390 ( .IN1(n1928), .IN2(n1929), .S(n2016), .Q(n1931) );
  NAND3X0 U2391 ( .IN1(\r[3][20] ), .IN2(n2015), .IN3(n2038), .QN(n1930) );
  MUX21X1 U2392 ( .IN1(n1932), .IN2(n1933), .S(n2016), .Q(n1935) );
  NAND3X0 U2393 ( .IN1(\r[3][19] ), .IN2(n2015), .IN3(n2038), .QN(n1934) );
  MUX21X1 U2394 ( .IN1(n1936), .IN2(n1937), .S(n2016), .Q(n1939) );
  NAND3X0 U2395 ( .IN1(\r[3][18] ), .IN2(n2015), .IN3(n2038), .QN(n1938) );
  MUX21X1 U2396 ( .IN1(n1940), .IN2(n1941), .S(n2016), .Q(n1943) );
  NAND3X0 U2397 ( .IN1(\r[3][17] ), .IN2(n2015), .IN3(n2038), .QN(n1942) );
  MUX21X1 U2398 ( .IN1(n1944), .IN2(n1945), .S(n2016), .Q(n1947) );
  NAND3X0 U2399 ( .IN1(\r[3][16] ), .IN2(n2015), .IN3(n2038), .QN(n1946) );
  MUX21X1 U2400 ( .IN1(n1948), .IN2(n1949), .S(n2016), .Q(n1951) );
  NAND3X0 U2401 ( .IN1(\r[3][15] ), .IN2(n2015), .IN3(n2038), .QN(n1950) );
  MUX21X1 U2402 ( .IN1(n1952), .IN2(n1953), .S(n2016), .Q(n1955) );
  NAND3X0 U2403 ( .IN1(\r[3][14] ), .IN2(n2015), .IN3(n2038), .QN(n1954) );
  MUX21X1 U2404 ( .IN1(n1956), .IN2(n1957), .S(n2016), .Q(n1959) );
  NAND3X0 U2405 ( .IN1(\r[3][13] ), .IN2(n2015), .IN3(n2038), .QN(n1958) );
  MUX21X1 U2406 ( .IN1(n1960), .IN2(n1961), .S(n2016), .Q(n1963) );
  NAND3X0 U2407 ( .IN1(\r[3][12] ), .IN2(n2014), .IN3(n2038), .QN(n1962) );
  MUX21X1 U2408 ( .IN1(n1964), .IN2(n1965), .S(n2016), .Q(n1967) );
  NAND3X0 U2409 ( .IN1(\r[3][11] ), .IN2(n2015), .IN3(n2038), .QN(n1966) );
  MUX21X1 U2410 ( .IN1(n1968), .IN2(n1969), .S(n2016), .Q(n1971) );
  NAND3X0 U2411 ( .IN1(\r[3][10] ), .IN2(n2014), .IN3(n2038), .QN(n1970) );
  MUX21X1 U2412 ( .IN1(n1972), .IN2(n1973), .S(n2016), .Q(n1975) );
  NAND3X0 U2413 ( .IN1(\r[3][9] ), .IN2(n2014), .IN3(n2038), .QN(n1974) );
  MUX21X1 U2414 ( .IN1(n1976), .IN2(n1977), .S(n2016), .Q(n1979) );
  NAND3X0 U2415 ( .IN1(\r[3][8] ), .IN2(n2014), .IN3(n2038), .QN(n1978) );
  MUX21X1 U2416 ( .IN1(n1980), .IN2(n1981), .S(n2016), .Q(n1983) );
  NAND3X0 U2417 ( .IN1(\r[3][7] ), .IN2(n2014), .IN3(n2038), .QN(n1982) );
  MUX21X1 U2418 ( .IN1(n1984), .IN2(n1985), .S(n2016), .Q(n1987) );
  NAND3X0 U2419 ( .IN1(\r[3][6] ), .IN2(n2014), .IN3(n2038), .QN(n1986) );
  MUX21X1 U2420 ( .IN1(n1988), .IN2(n1989), .S(n2016), .Q(n1991) );
  NAND3X0 U2421 ( .IN1(\r[3][5] ), .IN2(n2014), .IN3(n2038), .QN(n1990) );
  MUX21X1 U2422 ( .IN1(n1992), .IN2(n1993), .S(n2017), .Q(n1995) );
  NAND3X0 U2423 ( .IN1(\r[3][4] ), .IN2(n2014), .IN3(n2038), .QN(n1994) );
  MUX21X1 U2424 ( .IN1(n1996), .IN2(n1997), .S(n2017), .Q(n1999) );
  NAND3X0 U2425 ( .IN1(\r[3][3] ), .IN2(n2014), .IN3(n2038), .QN(n1998) );
  MUX21X1 U2426 ( .IN1(n2000), .IN2(n2001), .S(n2017), .Q(n2003) );
  NAND3X0 U2427 ( .IN1(\r[3][2] ), .IN2(n2014), .IN3(n2038), .QN(n2002) );
  MUX21X1 U2428 ( .IN1(n2004), .IN2(n2005), .S(n2017), .Q(n2007) );
  NAND3X0 U2429 ( .IN1(\r[3][1] ), .IN2(n2014), .IN3(n2038), .QN(n2006) );
  MUX21X1 U2430 ( .IN1(n2008), .IN2(n2009), .S(n2017), .Q(n2011) );
  NAND3X0 U2431 ( .IN1(\r[3][0] ), .IN2(n2015), .IN3(n2039), .QN(n2010) );
endmodule
